module hash_synth (target, clk, reset_L, num_entradas, bounty_synth_out, nonce_synth_valido_out, nonce_synth, fin_synth);

input clk;
input reset_L;
output fin_synth;
input [7:0] target;
input [1:0] num_entradas;
output [23:0] bounty_synth_out;
output [31:0] nonce_synth_valido_out;
output [31:0] nonce_synth;

wire vdd = 1'b1;
wire gnd = 1'b0;

	BUFX2 BUFX2_1 ( .A(clk), .Y(clk_hier0_bF_buf7) );
	BUFX2 BUFX2_2 ( .A(clk), .Y(clk_hier0_bF_buf6) );
	BUFX2 BUFX2_3 ( .A(clk), .Y(clk_hier0_bF_buf5) );
	BUFX2 BUFX2_4 ( .A(clk), .Y(clk_hier0_bF_buf4) );
	BUFX2 BUFX2_5 ( .A(clk), .Y(clk_hier0_bF_buf3) );
	BUFX2 BUFX2_6 ( .A(clk), .Y(clk_hier0_bF_buf2) );
	BUFX2 BUFX2_7 ( .A(clk), .Y(clk_hier0_bF_buf1) );
	BUFX2 BUFX2_8 ( .A(clk), .Y(clk_hier0_bF_buf0) );
	BUFX4 BUFX4_1 ( .A(_92_), .Y(_92__bF_buf6) );
	BUFX2 BUFX2_9 ( .A(_92_), .Y(_92__bF_buf5) );
	BUFX2 BUFX2_10 ( .A(_92_), .Y(_92__bF_buf4) );
	BUFX2 BUFX2_11 ( .A(_92_), .Y(_92__bF_buf3) );
	BUFX2 BUFX2_12 ( .A(_92_), .Y(_92__bF_buf2) );
	BUFX2 BUFX2_13 ( .A(_92_), .Y(_92__bF_buf1) );
	BUFX2 BUFX2_14 ( .A(_92_), .Y(_92__bF_buf0) );
	BUFX2 BUFX2_15 ( .A(_2633_), .Y(_2633__bF_buf6) );
	BUFX2 BUFX2_16 ( .A(_2633_), .Y(_2633__bF_buf5) );
	BUFX2 BUFX2_17 ( .A(_2633_), .Y(_2633__bF_buf4) );
	BUFX2 BUFX2_18 ( .A(_2633_), .Y(_2633__bF_buf3) );
	BUFX2 BUFX2_19 ( .A(_2633_), .Y(_2633__bF_buf2) );
	BUFX2 BUFX2_20 ( .A(_2633_), .Y(_2633__bF_buf1) );
	BUFX2 BUFX2_21 ( .A(_2633_), .Y(_2633__bF_buf0) );
	BUFX2 BUFX2_22 ( .A(_1202_), .Y(_1202__bF_buf5) );
	BUFX2 BUFX2_23 ( .A(_1202_), .Y(_1202__bF_buf4) );
	BUFX2 BUFX2_24 ( .A(_1202_), .Y(_1202__bF_buf3) );
	BUFX2 BUFX2_25 ( .A(_1202_), .Y(_1202__bF_buf2) );
	BUFX2 BUFX2_26 ( .A(_1202_), .Y(_1202__bF_buf1) );
	BUFX2 BUFX2_27 ( .A(_1202_), .Y(_1202__bF_buf0) );
	BUFX4 BUFX4_2 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf76) );
	BUFX4 BUFX4_3 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf75) );
	BUFX4 BUFX4_4 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf74) );
	BUFX4 BUFX4_5 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf73) );
	BUFX4 BUFX4_6 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf72) );
	BUFX4 BUFX4_7 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf71) );
	BUFX4 BUFX4_8 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf70) );
	BUFX4 BUFX4_9 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf69) );
	BUFX4 BUFX4_10 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf68) );
	BUFX4 BUFX4_11 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf67) );
	BUFX4 BUFX4_12 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf66) );
	BUFX4 BUFX4_13 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf65) );
	BUFX4 BUFX4_14 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf64) );
	BUFX4 BUFX4_15 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf63) );
	BUFX4 BUFX4_16 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf62) );
	BUFX4 BUFX4_17 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf61) );
	BUFX4 BUFX4_18 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf60) );
	BUFX4 BUFX4_19 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf59) );
	BUFX4 BUFX4_20 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf58) );
	BUFX4 BUFX4_21 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf57) );
	BUFX4 BUFX4_22 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf56) );
	BUFX4 BUFX4_23 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf55) );
	BUFX4 BUFX4_24 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf54) );
	BUFX4 BUFX4_25 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf53) );
	BUFX4 BUFX4_26 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf52) );
	BUFX4 BUFX4_27 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf51) );
	BUFX4 BUFX4_28 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf50) );
	BUFX4 BUFX4_29 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf49) );
	BUFX4 BUFX4_30 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf48) );
	BUFX4 BUFX4_31 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf47) );
	BUFX4 BUFX4_32 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf46) );
	BUFX4 BUFX4_33 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf45) );
	BUFX4 BUFX4_34 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf44) );
	BUFX4 BUFX4_35 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf43) );
	BUFX4 BUFX4_36 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf42) );
	BUFX4 BUFX4_37 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf41) );
	BUFX4 BUFX4_38 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf40) );
	BUFX4 BUFX4_39 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf39) );
	BUFX4 BUFX4_40 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf38) );
	BUFX4 BUFX4_41 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf37) );
	BUFX4 BUFX4_42 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf36) );
	BUFX4 BUFX4_43 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf35) );
	BUFX4 BUFX4_44 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf34) );
	BUFX4 BUFX4_45 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf33) );
	BUFX4 BUFX4_46 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf32) );
	BUFX4 BUFX4_47 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf31) );
	BUFX4 BUFX4_48 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf30) );
	BUFX4 BUFX4_49 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf29) );
	BUFX4 BUFX4_50 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf28) );
	BUFX4 BUFX4_51 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf27) );
	BUFX4 BUFX4_52 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf26) );
	BUFX4 BUFX4_53 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf25) );
	BUFX4 BUFX4_54 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf24) );
	BUFX4 BUFX4_55 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf23) );
	BUFX4 BUFX4_56 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf22) );
	BUFX4 BUFX4_57 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf21) );
	BUFX4 BUFX4_58 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf20) );
	BUFX4 BUFX4_59 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf19) );
	BUFX4 BUFX4_60 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf18) );
	BUFX4 BUFX4_61 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf17) );
	BUFX4 BUFX4_62 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf16) );
	BUFX4 BUFX4_63 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf15) );
	BUFX4 BUFX4_64 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf14) );
	BUFX4 BUFX4_65 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf13) );
	BUFX4 BUFX4_66 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf12) );
	BUFX4 BUFX4_67 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf11) );
	BUFX4 BUFX4_68 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf10) );
	BUFX4 BUFX4_69 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf9) );
	BUFX4 BUFX4_70 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf8) );
	BUFX4 BUFX4_71 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf7) );
	BUFX4 BUFX4_72 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf6) );
	BUFX4 BUFX4_73 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_74 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_75 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_76 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_77 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_78 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf0) );
	BUFX2 BUFX2_28 ( .A(_117_), .Y(_117__bF_buf6) );
	BUFX2 BUFX2_29 ( .A(_117_), .Y(_117__bF_buf5) );
	BUFX2 BUFX2_30 ( .A(_117_), .Y(_117__bF_buf4) );
	BUFX2 BUFX2_31 ( .A(_117_), .Y(_117__bF_buf3) );
	BUFX2 BUFX2_32 ( .A(_117_), .Y(_117__bF_buf2) );
	BUFX2 BUFX2_33 ( .A(_117_), .Y(_117__bF_buf1) );
	BUFX2 BUFX2_34 ( .A(_117_), .Y(_117__bF_buf0) );
	BUFX2 BUFX2_35 ( .A(_545_), .Y(_545__bF_buf4) );
	BUFX2 BUFX2_36 ( .A(_545_), .Y(_545__bF_buf3) );
	BUFX2 BUFX2_37 ( .A(_545_), .Y(_545__bF_buf2) );
	BUFX2 BUFX2_38 ( .A(_545_), .Y(_545__bF_buf1) );
	BUFX2 BUFX2_39 ( .A(_545_), .Y(_545__bF_buf0) );
	BUFX4 BUFX4_79 ( .A(_142_), .Y(_142__bF_buf6) );
	BUFX4 BUFX4_80 ( .A(_142_), .Y(_142__bF_buf5) );
	BUFX4 BUFX4_81 ( .A(_142_), .Y(_142__bF_buf4) );
	BUFX4 BUFX4_82 ( .A(_142_), .Y(_142__bF_buf3) );
	BUFX4 BUFX4_83 ( .A(_142_), .Y(_142__bF_buf2) );
	BUFX4 BUFX4_84 ( .A(_142_), .Y(_142__bF_buf1) );
	BUFX4 BUFX4_85 ( .A(_142_), .Y(_142__bF_buf0) );
	BUFX2 BUFX2_40 ( .A(_1549_), .Y(_1549__bF_buf3) );
	BUFX2 BUFX2_41 ( .A(_1549_), .Y(_1549__bF_buf2) );
	BUFX2 BUFX2_42 ( .A(_1549_), .Y(_1549__bF_buf1) );
	BUFX2 BUFX2_43 ( .A(_1549_), .Y(_1549__bF_buf0) );
	BUFX2 BUFX2_44 ( .A(_2470_), .Y(_2470__bF_buf3) );
	BUFX2 BUFX2_45 ( .A(_2470_), .Y(_2470__bF_buf2) );
	BUFX2 BUFX2_46 ( .A(_2470_), .Y(_2470__bF_buf1) );
	BUFX2 BUFX2_47 ( .A(_2470_), .Y(_2470__bF_buf0) );
	BUFX2 BUFX2_48 ( .A(_2625_), .Y(_2625__bF_buf6) );
	BUFX2 BUFX2_49 ( .A(_2625_), .Y(_2625__bF_buf5) );
	BUFX2 BUFX2_50 ( .A(_2625_), .Y(_2625__bF_buf4) );
	BUFX2 BUFX2_51 ( .A(_2625_), .Y(_2625__bF_buf3) );
	BUFX2 BUFX2_52 ( .A(_2625_), .Y(_2625__bF_buf2) );
	BUFX2 BUFX2_53 ( .A(_2625_), .Y(_2625__bF_buf1) );
	BUFX2 BUFX2_54 ( .A(_2625_), .Y(_2625__bF_buf0) );
	BUFX2 BUFX2_55 ( .A(_1379_), .Y(_1379__bF_buf3) );
	BUFX2 BUFX2_56 ( .A(_1379_), .Y(_1379__bF_buf2) );
	BUFX2 BUFX2_57 ( .A(_1379_), .Y(_1379__bF_buf1) );
	BUFX2 BUFX2_58 ( .A(_1379_), .Y(_1379__bF_buf0) );
	BUFX2 BUFX2_59 ( .A(_2618_), .Y(_2618__bF_buf6) );
	BUFX2 BUFX2_60 ( .A(_2618_), .Y(_2618__bF_buf5) );
	BUFX2 BUFX2_61 ( .A(_2618_), .Y(_2618__bF_buf4) );
	BUFX2 BUFX2_62 ( .A(_2618_), .Y(_2618__bF_buf3) );
	BUFX2 BUFX2_63 ( .A(_2618_), .Y(_2618__bF_buf2) );
	BUFX2 BUFX2_64 ( .A(_2618_), .Y(_2618__bF_buf1) );
	BUFX2 BUFX2_65 ( .A(_2618_), .Y(_2618__bF_buf0) );
	BUFX4 BUFX4_86 ( .A(_261_), .Y(_261__bF_buf15) );
	BUFX4 BUFX4_87 ( .A(_261_), .Y(_261__bF_buf14) );
	BUFX4 BUFX4_88 ( .A(_261_), .Y(_261__bF_buf13) );
	BUFX4 BUFX4_89 ( .A(_261_), .Y(_261__bF_buf12) );
	BUFX4 BUFX4_90 ( .A(_261_), .Y(_261__bF_buf11) );
	BUFX4 BUFX4_91 ( .A(_261_), .Y(_261__bF_buf10) );
	BUFX4 BUFX4_92 ( .A(_261_), .Y(_261__bF_buf9) );
	BUFX4 BUFX4_93 ( .A(_261_), .Y(_261__bF_buf8) );
	BUFX4 BUFX4_94 ( .A(_261_), .Y(_261__bF_buf7) );
	BUFX4 BUFX4_95 ( .A(_261_), .Y(_261__bF_buf6) );
	BUFX4 BUFX4_96 ( .A(_261_), .Y(_261__bF_buf5) );
	BUFX4 BUFX4_97 ( .A(_261_), .Y(_261__bF_buf4) );
	BUFX4 BUFX4_98 ( .A(_261_), .Y(_261__bF_buf3) );
	BUFX4 BUFX4_99 ( .A(_261_), .Y(_261__bF_buf2) );
	BUFX4 BUFX4_100 ( .A(_261_), .Y(_261__bF_buf1) );
	BUFX4 BUFX4_101 ( .A(_261_), .Y(_261__bF_buf0) );
	BUFX2 BUFX2_66 ( .A(_1205_), .Y(_1205__bF_buf3) );
	BUFX2 BUFX2_67 ( .A(_1205_), .Y(_1205__bF_buf2) );
	BUFX2 BUFX2_68 ( .A(_1205_), .Y(_1205__bF_buf1) );
	BUFX2 BUFX2_69 ( .A(_1205_), .Y(_1205__bF_buf0) );
	BUFX2 BUFX2_70 ( .A(_53_), .Y(_53__bF_buf6) );
	BUFX2 BUFX2_71 ( .A(_53_), .Y(_53__bF_buf5) );
	BUFX2 BUFX2_72 ( .A(_53_), .Y(_53__bF_buf4) );
	BUFX2 BUFX2_73 ( .A(_53_), .Y(_53__bF_buf3) );
	BUFX2 BUFX2_74 ( .A(_53_), .Y(_53__bF_buf2) );
	BUFX2 BUFX2_75 ( .A(_53_), .Y(_53__bF_buf1) );
	BUFX2 BUFX2_76 ( .A(_53_), .Y(_53__bF_buf0) );
	BUFX2 BUFX2_77 ( .A(_2189_), .Y(_2189__bF_buf4) );
	BUFX2 BUFX2_78 ( .A(_2189_), .Y(_2189__bF_buf3) );
	BUFX2 BUFX2_79 ( .A(_2189_), .Y(_2189__bF_buf2) );
	BUFX2 BUFX2_80 ( .A(_2189_), .Y(_2189__bF_buf1) );
	BUFX2 BUFX2_81 ( .A(_2189_), .Y(_2189__bF_buf0) );
	BUFX2 BUFX2_82 ( .A(comparador_valid), .Y(comparador_valid_bF_buf5) );
	BUFX4 BUFX4_102 ( .A(comparador_valid), .Y(comparador_valid_bF_buf4) );
	BUFX2 BUFX2_83 ( .A(comparador_valid), .Y(comparador_valid_bF_buf3) );
	BUFX2 BUFX2_84 ( .A(comparador_valid), .Y(comparador_valid_bF_buf2) );
	BUFX2 BUFX2_85 ( .A(comparador_valid), .Y(comparador_valid_bF_buf1) );
	BUFX2 BUFX2_86 ( .A(comparador_valid), .Y(comparador_valid_bF_buf0) );
	BUFX2 BUFX2_87 ( .A(_1380_), .Y(_1380__bF_buf6) );
	BUFX2 BUFX2_88 ( .A(_1380_), .Y(_1380__bF_buf5) );
	BUFX2 BUFX2_89 ( .A(_1380_), .Y(_1380__bF_buf4) );
	BUFX2 BUFX2_90 ( .A(_1380_), .Y(_1380__bF_buf3) );
	BUFX2 BUFX2_91 ( .A(_1380_), .Y(_1380__bF_buf2) );
	BUFX2 BUFX2_92 ( .A(_1380_), .Y(_1380__bF_buf1) );
	BUFX2 BUFX2_93 ( .A(_1380_), .Y(_1380__bF_buf0) );
	BUFX2 BUFX2_94 ( .A(_1547_), .Y(_1547__bF_buf3) );
	BUFX2 BUFX2_95 ( .A(_1547_), .Y(_1547__bF_buf2) );
	BUFX2 BUFX2_96 ( .A(_1547_), .Y(_1547__bF_buf1) );
	BUFX2 BUFX2_97 ( .A(_1547_), .Y(_1547__bF_buf0) );
	BUFX4 BUFX4_103 ( .A(_2473_), .Y(_2473__bF_buf15) );
	BUFX4 BUFX4_104 ( .A(_2473_), .Y(_2473__bF_buf14) );
	BUFX4 BUFX4_105 ( .A(_2473_), .Y(_2473__bF_buf13) );
	BUFX4 BUFX4_106 ( .A(_2473_), .Y(_2473__bF_buf12) );
	BUFX4 BUFX4_107 ( .A(_2473_), .Y(_2473__bF_buf11) );
	BUFX4 BUFX4_108 ( .A(_2473_), .Y(_2473__bF_buf10) );
	BUFX4 BUFX4_109 ( .A(_2473_), .Y(_2473__bF_buf9) );
	BUFX4 BUFX4_110 ( .A(_2473_), .Y(_2473__bF_buf8) );
	BUFX4 BUFX4_111 ( .A(_2473_), .Y(_2473__bF_buf7) );
	BUFX4 BUFX4_112 ( .A(_2473_), .Y(_2473__bF_buf6) );
	BUFX4 BUFX4_113 ( .A(_2473_), .Y(_2473__bF_buf5) );
	BUFX4 BUFX4_114 ( .A(_2473_), .Y(_2473__bF_buf4) );
	BUFX4 BUFX4_115 ( .A(_2473_), .Y(_2473__bF_buf3) );
	BUFX4 BUFX4_116 ( .A(_2473_), .Y(_2473__bF_buf2) );
	BUFX4 BUFX4_117 ( .A(_2473_), .Y(_2473__bF_buf1) );
	BUFX4 BUFX4_118 ( .A(_2473_), .Y(_2473__bF_buf0) );
	BUFX2 BUFX2_98 ( .A(_1373_), .Y(_1373__bF_buf3) );
	BUFX2 BUFX2_99 ( .A(_1373_), .Y(_1373__bF_buf2) );
	BUFX2 BUFX2_100 ( .A(_1373_), .Y(_1373__bF_buf1) );
	BUFX2 BUFX2_101 ( .A(_1373_), .Y(_1373__bF_buf0) );
	BUFX2 BUFX2_102 ( .A(_1269_), .Y(_1269__bF_buf3) );
	BUFX2 BUFX2_103 ( .A(_1269_), .Y(_1269__bF_buf2) );
	BUFX2 BUFX2_104 ( .A(_1269_), .Y(_1269__bF_buf1) );
	BUFX2 BUFX2_105 ( .A(_1269_), .Y(_1269__bF_buf0) );
	BUFX4 BUFX4_119 ( .A(concatenador_count_1_), .Y(concatenador_count_1_bF_buf6) );
	BUFX4 BUFX4_120 ( .A(concatenador_count_1_), .Y(concatenador_count_1_bF_buf5) );
	BUFX4 BUFX4_121 ( .A(concatenador_count_1_), .Y(concatenador_count_1_bF_buf4) );
	BUFX4 BUFX4_122 ( .A(concatenador_count_1_), .Y(concatenador_count_1_bF_buf3) );
	BUFX4 BUFX4_123 ( .A(concatenador_count_1_), .Y(concatenador_count_1_bF_buf2) );
	BUFX4 BUFX4_124 ( .A(concatenador_count_1_), .Y(concatenador_count_1_bF_buf1) );
	BUFX4 BUFX4_125 ( .A(concatenador_count_1_), .Y(concatenador_count_1_bF_buf0) );
	BUFX2 BUFX2_106 ( .A(_1354_), .Y(_1354__bF_buf3) );
	BUFX2 BUFX2_107 ( .A(_1354_), .Y(_1354__bF_buf2) );
	BUFX2 BUFX2_108 ( .A(_1354_), .Y(_1354__bF_buf1) );
	BUFX2 BUFX2_109 ( .A(_1354_), .Y(_1354__bF_buf0) );
	BUFX2 BUFX2_110 ( .A(_10_), .Y(_10__bF_buf6) );
	BUFX2 BUFX2_111 ( .A(_10_), .Y(_10__bF_buf5) );
	BUFX2 BUFX2_112 ( .A(_10_), .Y(_10__bF_buf4) );
	BUFX2 BUFX2_113 ( .A(_10_), .Y(_10__bF_buf3) );
	BUFX2 BUFX2_114 ( .A(_10_), .Y(_10__bF_buf2) );
	BUFX2 BUFX2_115 ( .A(_10_), .Y(_10__bF_buf1) );
	BUFX2 BUFX2_116 ( .A(_10_), .Y(_10__bF_buf0) );
	BUFX2 BUFX2_117 ( .A(_1_), .Y(_1__bF_buf5) );
	BUFX2 BUFX2_118 ( .A(_1_), .Y(_1__bF_buf4) );
	BUFX2 BUFX2_119 ( .A(_1_), .Y(_1__bF_buf3) );
	BUFX2 BUFX2_120 ( .A(_1_), .Y(_1__bF_buf2) );
	BUFX2 BUFX2_121 ( .A(_1_), .Y(_1__bF_buf1) );
	BUFX2 BUFX2_122 ( .A(_1_), .Y(_1__bF_buf0) );
	BUFX4 BUFX4_126 ( .A(reset_L), .Y(reset_L_bF_buf11) );
	BUFX4 BUFX4_127 ( .A(reset_L), .Y(reset_L_bF_buf10) );
	BUFX4 BUFX4_128 ( .A(reset_L), .Y(reset_L_bF_buf9) );
	BUFX4 BUFX4_129 ( .A(reset_L), .Y(reset_L_bF_buf8) );
	BUFX4 BUFX4_130 ( .A(reset_L), .Y(reset_L_bF_buf7) );
	BUFX4 BUFX4_131 ( .A(reset_L), .Y(reset_L_bF_buf6) );
	BUFX4 BUFX4_132 ( .A(reset_L), .Y(reset_L_bF_buf5) );
	BUFX4 BUFX4_133 ( .A(reset_L), .Y(reset_L_bF_buf4) );
	BUFX4 BUFX4_134 ( .A(reset_L), .Y(reset_L_bF_buf3) );
	BUFX4 BUFX4_135 ( .A(reset_L), .Y(reset_L_bF_buf2) );
	BUFX4 BUFX4_136 ( .A(reset_L), .Y(reset_L_bF_buf1) );
	BUFX4 BUFX4_137 ( .A(reset_L), .Y(reset_L_bF_buf0) );
	BUFX2 BUFX2_123 ( .A(_558_), .Y(_558__bF_buf3) );
	BUFX2 BUFX2_124 ( .A(_558_), .Y(_558__bF_buf2) );
	BUFX2 BUFX2_125 ( .A(_558_), .Y(_558__bF_buf1) );
	BUFX2 BUFX2_126 ( .A(_558_), .Y(_558__bF_buf0) );
	BUFX2 BUFX2_127 ( .A(_2609_), .Y(_2609__bF_buf3) );
	BUFX2 BUFX2_128 ( .A(_2609_), .Y(_2609__bF_buf2) );
	BUFX2 BUFX2_129 ( .A(_2609_), .Y(_2609__bF_buf1) );
	BUFX2 BUFX2_130 ( .A(_2609_), .Y(_2609__bF_buf0) );
	BUFX2 BUFX2_131 ( .A(_1196_), .Y(_1196__bF_buf3) );
	BUFX2 BUFX2_132 ( .A(_1196_), .Y(_1196__bF_buf2) );
	BUFX2 BUFX2_133 ( .A(_1196_), .Y(_1196__bF_buf1) );
	BUFX2 BUFX2_134 ( .A(_1196_), .Y(_1196__bF_buf0) );
	BUFX4 BUFX4_138 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf11) );
	BUFX4 BUFX4_139 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf10) );
	BUFX4 BUFX4_140 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf9) );
	BUFX4 BUFX4_141 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf8) );
	BUFX4 BUFX4_142 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf7) );
	BUFX4 BUFX4_143 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf6) );
	BUFX4 BUFX4_144 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf5) );
	BUFX4 BUFX4_145 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf4) );
	BUFX4 BUFX4_146 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf3) );
	BUFX4 BUFX4_147 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf2) );
	BUFX4 BUFX4_148 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf1) );
	BUFX4 BUFX4_149 ( .A(concatenador_count_0_), .Y(concatenador_count_0_bF_buf0) );
	BUFX4 BUFX4_150 ( .A(_2471_), .Y(_2471__bF_buf13) );
	BUFX4 BUFX4_151 ( .A(_2471_), .Y(_2471__bF_buf12) );
	BUFX4 BUFX4_152 ( .A(_2471_), .Y(_2471__bF_buf11) );
	BUFX4 BUFX4_153 ( .A(_2471_), .Y(_2471__bF_buf10) );
	BUFX4 BUFX4_154 ( .A(_2471_), .Y(_2471__bF_buf9) );
	BUFX4 BUFX4_155 ( .A(_2471_), .Y(_2471__bF_buf8) );
	BUFX4 BUFX4_156 ( .A(_2471_), .Y(_2471__bF_buf7) );
	BUFX4 BUFX4_157 ( .A(_2471_), .Y(_2471__bF_buf6) );
	BUFX4 BUFX4_158 ( .A(_2471_), .Y(_2471__bF_buf5) );
	BUFX4 BUFX4_159 ( .A(_2471_), .Y(_2471__bF_buf4) );
	BUFX4 BUFX4_160 ( .A(_2471_), .Y(_2471__bF_buf3) );
	BUFX4 BUFX4_161 ( .A(_2471_), .Y(_2471__bF_buf2) );
	BUFX4 BUFX4_162 ( .A(_2471_), .Y(_2471__bF_buf1) );
	BUFX4 BUFX4_163 ( .A(_2471_), .Y(_2471__bF_buf0) );
	BUFX2 BUFX2_135 ( .A(_0__0_), .Y(bounty_synth_out[0]) );
	BUFX2 BUFX2_136 ( .A(_0__1_), .Y(bounty_synth_out[1]) );
	BUFX2 BUFX2_137 ( .A(_0__2_), .Y(bounty_synth_out[2]) );
	BUFX2 BUFX2_138 ( .A(_0__3_), .Y(bounty_synth_out[3]) );
	BUFX2 BUFX2_139 ( .A(_0__4_), .Y(bounty_synth_out[4]) );
	BUFX2 BUFX2_140 ( .A(_0__5_), .Y(bounty_synth_out[5]) );
	BUFX2 BUFX2_141 ( .A(_0__6_), .Y(bounty_synth_out[6]) );
	BUFX2 BUFX2_142 ( .A(_0__7_), .Y(bounty_synth_out[7]) );
	BUFX2 BUFX2_143 ( .A(_0__8_), .Y(bounty_synth_out[8]) );
	BUFX2 BUFX2_144 ( .A(_0__9_), .Y(bounty_synth_out[9]) );
	BUFX2 BUFX2_145 ( .A(_0__10_), .Y(bounty_synth_out[10]) );
	BUFX2 BUFX2_146 ( .A(_0__11_), .Y(bounty_synth_out[11]) );
	BUFX2 BUFX2_147 ( .A(_0__12_), .Y(bounty_synth_out[12]) );
	BUFX2 BUFX2_148 ( .A(_0__13_), .Y(bounty_synth_out[13]) );
	BUFX2 BUFX2_149 ( .A(_0__14_), .Y(bounty_synth_out[14]) );
	BUFX2 BUFX2_150 ( .A(_0__15_), .Y(bounty_synth_out[15]) );
	BUFX2 BUFX2_151 ( .A(_0__16_), .Y(bounty_synth_out[16]) );
	BUFX2 BUFX2_152 ( .A(_0__17_), .Y(bounty_synth_out[17]) );
	BUFX2 BUFX2_153 ( .A(_0__18_), .Y(bounty_synth_out[18]) );
	BUFX2 BUFX2_154 ( .A(_0__19_), .Y(bounty_synth_out[19]) );
	BUFX2 BUFX2_155 ( .A(_0__20_), .Y(bounty_synth_out[20]) );
	BUFX2 BUFX2_156 ( .A(_0__21_), .Y(bounty_synth_out[21]) );
	BUFX2 BUFX2_157 ( .A(_0__22_), .Y(bounty_synth_out[22]) );
	BUFX2 BUFX2_158 ( .A(_0__23_), .Y(bounty_synth_out[23]) );
	BUFX2 BUFX2_159 ( .A(_1__bF_buf5), .Y(fin_synth) );
	BUFX2 BUFX2_160 ( .A(_2__0_), .Y(nonce_synth[0]) );
	BUFX2 BUFX2_161 ( .A(_2__1_), .Y(nonce_synth[1]) );
	BUFX2 BUFX2_162 ( .A(_2__2_), .Y(nonce_synth[2]) );
	BUFX2 BUFX2_163 ( .A(_2__3_), .Y(nonce_synth[3]) );
	BUFX2 BUFX2_164 ( .A(_2__4_), .Y(nonce_synth[4]) );
	BUFX2 BUFX2_165 ( .A(_2__5_), .Y(nonce_synth[5]) );
	BUFX2 BUFX2_166 ( .A(_2__6_), .Y(nonce_synth[6]) );
	BUFX2 BUFX2_167 ( .A(_2__7_), .Y(nonce_synth[7]) );
	BUFX2 BUFX2_168 ( .A(_2__8_), .Y(nonce_synth[8]) );
	BUFX2 BUFX2_169 ( .A(_2__9_), .Y(nonce_synth[9]) );
	BUFX2 BUFX2_170 ( .A(_2__10_), .Y(nonce_synth[10]) );
	BUFX2 BUFX2_171 ( .A(_2__11_), .Y(nonce_synth[11]) );
	BUFX2 BUFX2_172 ( .A(_2__12_), .Y(nonce_synth[12]) );
	BUFX2 BUFX2_173 ( .A(_2__13_), .Y(nonce_synth[13]) );
	BUFX2 BUFX2_174 ( .A(_2__14_), .Y(nonce_synth[14]) );
	BUFX2 BUFX2_175 ( .A(_2__15_), .Y(nonce_synth[15]) );
	BUFX2 BUFX2_176 ( .A(_2__16_), .Y(nonce_synth[16]) );
	BUFX2 BUFX2_177 ( .A(_2__17_), .Y(nonce_synth[17]) );
	BUFX2 BUFX2_178 ( .A(_2__18_), .Y(nonce_synth[18]) );
	BUFX2 BUFX2_179 ( .A(_2__19_), .Y(nonce_synth[19]) );
	BUFX2 BUFX2_180 ( .A(_2__20_), .Y(nonce_synth[20]) );
	BUFX2 BUFX2_181 ( .A(_2__21_), .Y(nonce_synth[21]) );
	BUFX2 BUFX2_182 ( .A(_2__22_), .Y(nonce_synth[22]) );
	BUFX2 BUFX2_183 ( .A(_2__23_), .Y(nonce_synth[23]) );
	BUFX2 BUFX2_184 ( .A(_2__24_), .Y(nonce_synth[24]) );
	BUFX2 BUFX2_185 ( .A(_2__25_), .Y(nonce_synth[25]) );
	BUFX2 BUFX2_186 ( .A(_2__26_), .Y(nonce_synth[26]) );
	BUFX2 BUFX2_187 ( .A(_2__27_), .Y(nonce_synth[27]) );
	BUFX2 BUFX2_188 ( .A(_2__28_), .Y(nonce_synth[28]) );
	BUFX2 BUFX2_189 ( .A(_2__29_), .Y(nonce_synth[29]) );
	BUFX2 BUFX2_190 ( .A(_2__30_), .Y(nonce_synth[30]) );
	BUFX2 BUFX2_191 ( .A(_2__31_), .Y(nonce_synth[31]) );
	BUFX2 BUFX2_192 ( .A(_3__0_), .Y(nonce_synth_valido_out[0]) );
	BUFX2 BUFX2_193 ( .A(_3__1_), .Y(nonce_synth_valido_out[1]) );
	BUFX2 BUFX2_194 ( .A(_3__2_), .Y(nonce_synth_valido_out[2]) );
	BUFX2 BUFX2_195 ( .A(_3__3_), .Y(nonce_synth_valido_out[3]) );
	BUFX2 BUFX2_196 ( .A(_3__4_), .Y(nonce_synth_valido_out[4]) );
	BUFX2 BUFX2_197 ( .A(_3__5_), .Y(nonce_synth_valido_out[5]) );
	BUFX2 BUFX2_198 ( .A(_3__6_), .Y(nonce_synth_valido_out[6]) );
	BUFX2 BUFX2_199 ( .A(_3__7_), .Y(nonce_synth_valido_out[7]) );
	BUFX2 BUFX2_200 ( .A(_3__8_), .Y(nonce_synth_valido_out[8]) );
	BUFX2 BUFX2_201 ( .A(_3__9_), .Y(nonce_synth_valido_out[9]) );
	BUFX2 BUFX2_202 ( .A(_3__10_), .Y(nonce_synth_valido_out[10]) );
	BUFX2 BUFX2_203 ( .A(_3__11_), .Y(nonce_synth_valido_out[11]) );
	BUFX2 BUFX2_204 ( .A(_3__12_), .Y(nonce_synth_valido_out[12]) );
	BUFX2 BUFX2_205 ( .A(_3__13_), .Y(nonce_synth_valido_out[13]) );
	BUFX2 BUFX2_206 ( .A(_3__14_), .Y(nonce_synth_valido_out[14]) );
	BUFX2 BUFX2_207 ( .A(_3__15_), .Y(nonce_synth_valido_out[15]) );
	BUFX2 BUFX2_208 ( .A(_3__16_), .Y(nonce_synth_valido_out[16]) );
	BUFX2 BUFX2_209 ( .A(_3__17_), .Y(nonce_synth_valido_out[17]) );
	BUFX2 BUFX2_210 ( .A(_3__18_), .Y(nonce_synth_valido_out[18]) );
	BUFX2 BUFX2_211 ( .A(_3__19_), .Y(nonce_synth_valido_out[19]) );
	BUFX2 BUFX2_212 ( .A(_3__20_), .Y(nonce_synth_valido_out[20]) );
	BUFX2 BUFX2_213 ( .A(_3__21_), .Y(nonce_synth_valido_out[21]) );
	BUFX2 BUFX2_214 ( .A(_3__22_), .Y(nonce_synth_valido_out[22]) );
	BUFX2 BUFX2_215 ( .A(_3__23_), .Y(nonce_synth_valido_out[23]) );
	BUFX2 BUFX2_216 ( .A(_3__24_), .Y(nonce_synth_valido_out[24]) );
	BUFX2 BUFX2_217 ( .A(_3__25_), .Y(nonce_synth_valido_out[25]) );
	BUFX2 BUFX2_218 ( .A(_3__26_), .Y(nonce_synth_valido_out[26]) );
	BUFX2 BUFX2_219 ( .A(_3__27_), .Y(nonce_synth_valido_out[27]) );
	BUFX2 BUFX2_220 ( .A(_3__28_), .Y(nonce_synth_valido_out[28]) );
	BUFX2 BUFX2_221 ( .A(_3__29_), .Y(nonce_synth_valido_out[29]) );
	BUFX2 BUFX2_222 ( .A(_3__30_), .Y(nonce_synth_valido_out[30]) );
	BUFX2 BUFX2_223 ( .A(_3__31_), .Y(nonce_synth_valido_out[31]) );
	NAND2X1 NAND2X1_1 ( .A(reset_L_bF_buf11), .B(RAM_rd_ptr_0_), .Y(_4__88_) );
	INVX1 INVX1_1 ( .A(_4__88_), .Y(_4__89_) );
	NAND2X1 NAND2X1_2 ( .A(reset_L_bF_buf10), .B(RAM_rd_ptr_1_), .Y(_4__92_) );
	INVX1 INVX1_2 ( .A(_4__92_), .Y(_4__77_) );
	OR2X2 OR2X2_1 ( .A(_4__88_), .B(RAM_rd_ptr_1_), .Y(_4__84_) );
	NOR2X1 NOR2X1_1 ( .A(RAM_rd_ptr_0_), .B(_4__92_), .Y(_4__94_) );
	NAND3X1 NAND3X1_1 ( .A(reset_L_bF_buf9), .B(RAM_rd_ptr_0_), .C(RAM_rd_ptr_1_), .Y(_4__93_) );
	OAI21X1 OAI21X1_1 ( .A(RAM_rd_ptr_0_), .B(RAM_rd_ptr_1_), .C(reset_L_bF_buf8), .Y(_4__82_) );
	INVX1 INVX1_3 ( .A(_4__82_), .Y(_4__95_) );
	NAND2X1 NAND2X1_3 ( .A(RAM_rd_ptr_0_), .B(RAM_rd_ptr_1_), .Y(_5_) );
	OR2X2 OR2X2_2 ( .A(RAM_rd_ptr_0_), .B(RAM_rd_ptr_1_), .Y(_6_) );
	NAND3X1 NAND3X1_2 ( .A(reset_L_bF_buf7), .B(_5_), .C(_6_), .Y(_4__86_) );
	AOI21X1 AOI21X1_1 ( .A(RAM_rd_ptr_0_), .B(RAM_rd_ptr_1_), .C(_4__82_), .Y(_4__46_) );
	INVX1 INVX1_4 ( .A(_4__93_), .Y(_4__71_) );
	NOR2X1 NOR2X1_2 ( .A(RAM_rd_ptr_1_), .B(_4__88_), .Y(_4__58_) );
	OR2X2 OR2X2_3 ( .A(_4__92_), .B(RAM_rd_ptr_0_), .Y(_4__85_) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf76), .D(_4__46_), .Q(RAM_entrada_46_) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf75), .D(_4__58_), .Q(RAM_entrada_58_) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf74), .D(_4__95_), .Q(RAM_entrada_95_) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf73), .D(_4__71_), .Q(RAM_entrada_71_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf72), .D(_4__77_), .Q(RAM_entrada_77_) );
	DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf71), .D(_4__82_), .Q(RAM_entrada_82_) );
	DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf70), .D(_4__84_), .Q(RAM_entrada_84_) );
	DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf69), .D(_4__85_), .Q(RAM_entrada_85_) );
	DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf68), .D(_4__86_), .Q(RAM_entrada_86_) );
	DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf67), .D(_4__88_), .Q(RAM_entrada_88_) );
	DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf66), .D(_4__89_), .Q(RAM_entrada_89_) );
	DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf65), .D(_4__92_), .Q(RAM_entrada_92_) );
	DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf64), .D(_4__93_), .Q(RAM_entrada_93_) );
	DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf63), .D(_4__94_), .Q(RAM_entrada_94_) );
	INVX8 INVX8_1 ( .A(reset_L_bF_buf6), .Y(_10_) );
	INVX1 INVX1_5 ( .A(H_17_), .Y(_11_) );
	NOR2X1 NOR2X1_3 ( .A(target[1]), .B(_11_), .Y(_12_) );
	INVX1 INVX1_6 ( .A(H_16_), .Y(_13_) );
	NAND2X1 NAND2X1_4 ( .A(target[0]), .B(_13_), .Y(_14_) );
	NAND2X1 NAND2X1_5 ( .A(target[1]), .B(_11_), .Y(_15_) );
	AOI21X1 AOI21X1_2 ( .A(_14_), .B(_15_), .C(_12_), .Y(_16_) );
	AND2X2 AND2X2_1 ( .A(target[3]), .B(H_19_), .Y(_17_) );
	NOR2X1 NOR2X1_4 ( .A(target[3]), .B(H_19_), .Y(_18_) );
	NAND2X1 NAND2X1_6 ( .A(target[2]), .B(H_18_), .Y(_19_) );
	INVX1 INVX1_7 ( .A(_19_), .Y(_20_) );
	NOR2X1 NOR2X1_5 ( .A(target[2]), .B(H_18_), .Y(_21_) );
	OAI22X1 OAI22X1_1 ( .A(_17_), .B(_18_), .C(_20_), .D(_21_), .Y(_22_) );
	INVX1 INVX1_8 ( .A(H_19_), .Y(_23_) );
	NOR2X1 NOR2X1_6 ( .A(target[3]), .B(_23_), .Y(_24_) );
	NAND2X1 NAND2X1_7 ( .A(target[3]), .B(_23_), .Y(_25_) );
	INVX1 INVX1_9 ( .A(H_18_), .Y(_26_) );
	NOR2X1 NOR2X1_7 ( .A(target[2]), .B(_26_), .Y(_27_) );
	AOI21X1 AOI21X1_3 ( .A(_25_), .B(_27_), .C(_24_), .Y(_28_) );
	OAI21X1 OAI21X1_2 ( .A(_22_), .B(_16_), .C(_28_), .Y(_29_) );
	NAND2X1 NAND2X1_8 ( .A(target[7]), .B(H_23_), .Y(_30_) );
	INVX1 INVX1_10 ( .A(_30_), .Y(_31_) );
	NOR2X1 NOR2X1_8 ( .A(target[7]), .B(H_23_), .Y(_32_) );
	NAND2X1 NAND2X1_9 ( .A(target[6]), .B(H_22_), .Y(_33_) );
	INVX1 INVX1_11 ( .A(_33_), .Y(_34_) );
	NOR2X1 NOR2X1_9 ( .A(target[6]), .B(H_22_), .Y(_35_) );
	OAI22X1 OAI22X1_2 ( .A(_31_), .B(_32_), .C(_34_), .D(_35_), .Y(_36_) );
	INVX1 INVX1_12 ( .A(target[5]), .Y(_37_) );
	INVX1 INVX1_13 ( .A(target[4]), .Y(_38_) );
	AOI22X1 AOI22X1_1 ( .A(_37_), .B(H_21_), .C(_38_), .D(H_20_), .Y(_39_) );
	INVX1 INVX1_14 ( .A(H_21_), .Y(_40_) );
	INVX1 INVX1_15 ( .A(H_20_), .Y(_41_) );
	AOI22X1 AOI22X1_2 ( .A(_40_), .B(target[5]), .C(target[4]), .D(_41_), .Y(_42_) );
	NAND2X1 NAND2X1_10 ( .A(_39_), .B(_42_), .Y(_43_) );
	NOR2X1 NOR2X1_10 ( .A(_36_), .B(_43_), .Y(_44_) );
	INVX1 INVX1_16 ( .A(target[7]), .Y(_45_) );
	INVX1 INVX1_17 ( .A(H_23_), .Y(_46_) );
	INVX1 INVX1_18 ( .A(H_22_), .Y(_47_) );
	OAI22X1 OAI22X1_3 ( .A(_46_), .B(target[7]), .C(target[6]), .D(_47_), .Y(_48_) );
	OAI21X1 OAI21X1_3 ( .A(_45_), .B(H_23_), .C(_48_), .Y(_49_) );
	OAI22X1 OAI22X1_4 ( .A(_40_), .B(target[5]), .C(target[4]), .D(_41_), .Y(_50_) );
	OAI21X1 OAI21X1_4 ( .A(_37_), .B(H_21_), .C(_50_), .Y(_51_) );
	OAI21X1 OAI21X1_5 ( .A(_51_), .B(_36_), .C(_49_), .Y(_52_) );
	AOI21X1 AOI21X1_4 ( .A(_44_), .B(_29_), .C(_52_), .Y(_53_) );
	INVX1 INVX1_19 ( .A(H_9_), .Y(_54_) );
	NOR2X1 NOR2X1_11 ( .A(target[1]), .B(_54_), .Y(_55_) );
	INVX1 INVX1_20 ( .A(H_8_), .Y(_56_) );
	NAND2X1 NAND2X1_11 ( .A(target[0]), .B(_56_), .Y(_57_) );
	NAND2X1 NAND2X1_12 ( .A(target[1]), .B(_54_), .Y(_58_) );
	AOI21X1 AOI21X1_5 ( .A(_57_), .B(_58_), .C(_55_), .Y(_59_) );
	NAND2X1 NAND2X1_13 ( .A(target[3]), .B(H_11_), .Y(_60_) );
	INVX1 INVX1_21 ( .A(_60_), .Y(_61_) );
	NOR2X1 NOR2X1_12 ( .A(target[3]), .B(H_11_), .Y(_62_) );
	NAND2X1 NAND2X1_14 ( .A(target[2]), .B(H_10_), .Y(_63_) );
	INVX1 INVX1_22 ( .A(_63_), .Y(_64_) );
	NOR2X1 NOR2X1_13 ( .A(target[2]), .B(H_10_), .Y(_65_) );
	OAI22X1 OAI22X1_5 ( .A(_61_), .B(_62_), .C(_64_), .D(_65_), .Y(_66_) );
	INVX1 INVX1_23 ( .A(H_11_), .Y(_67_) );
	NOR2X1 NOR2X1_14 ( .A(target[3]), .B(_67_), .Y(_68_) );
	NAND2X1 NAND2X1_15 ( .A(target[3]), .B(_67_), .Y(_69_) );
	INVX1 INVX1_24 ( .A(H_10_), .Y(_70_) );
	NOR2X1 NOR2X1_15 ( .A(target[2]), .B(_70_), .Y(_71_) );
	AOI21X1 AOI21X1_6 ( .A(_69_), .B(_71_), .C(_68_), .Y(_72_) );
	OAI21X1 OAI21X1_6 ( .A(_66_), .B(_59_), .C(_72_), .Y(_73_) );
	INVX1 INVX1_25 ( .A(H_14_), .Y(_74_) );
	NAND2X1 NAND2X1_16 ( .A(target[6]), .B(_74_), .Y(_75_) );
	INVX1 INVX1_26 ( .A(H_15_), .Y(_76_) );
	NAND2X1 NAND2X1_17 ( .A(target[7]), .B(_76_), .Y(_77_) );
	INVX1 INVX1_27 ( .A(target[6]), .Y(_78_) );
	AOI22X1 AOI22X1_3 ( .A(_45_), .B(H_15_), .C(_78_), .D(H_14_), .Y(_79_) );
	NAND3X1 NAND3X1_3 ( .A(_75_), .B(_77_), .C(_79_), .Y(_80_) );
	AOI22X1 AOI22X1_4 ( .A(_37_), .B(H_13_), .C(_38_), .D(H_12_), .Y(_81_) );
	INVX1 INVX1_28 ( .A(H_13_), .Y(_82_) );
	INVX1 INVX1_29 ( .A(H_12_), .Y(_83_) );
	AOI22X1 AOI22X1_5 ( .A(_82_), .B(target[5]), .C(target[4]), .D(_83_), .Y(_84_) );
	NAND2X1 NAND2X1_18 ( .A(_81_), .B(_84_), .Y(_85_) );
	NOR2X1 NOR2X1_16 ( .A(_85_), .B(_80_), .Y(_86_) );
	OAI22X1 OAI22X1_6 ( .A(_82_), .B(target[5]), .C(target[4]), .D(_83_), .Y(_87_) );
	OAI21X1 OAI21X1_7 ( .A(_37_), .B(H_13_), .C(_87_), .Y(_88_) );
	OAI22X1 OAI22X1_7 ( .A(_76_), .B(target[7]), .C(target[6]), .D(_74_), .Y(_89_) );
	AOI21X1 AOI21X1_7 ( .A(_77_), .B(_89_), .C(_1__bF_buf4), .Y(_90_) );
	OAI21X1 OAI21X1_8 ( .A(_80_), .B(_88_), .C(_90_), .Y(_91_) );
	AOI21X1 AOI21X1_8 ( .A(_73_), .B(_86_), .C(_91_), .Y(_92_) );
	NAND3X1 NAND3X1_4 ( .A(H_0_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_93_) );
	INVX1 INVX1_30 ( .A(target[1]), .Y(_94_) );
	NAND2X1 NAND2X1_19 ( .A(H_17_), .B(_94_), .Y(_95_) );
	INVX1 INVX1_31 ( .A(target[0]), .Y(_96_) );
	OAI22X1 OAI22X1_8 ( .A(_94_), .B(H_17_), .C(_96_), .D(H_16_), .Y(_97_) );
	NAND2X1 NAND2X1_20 ( .A(_95_), .B(_97_), .Y(_98_) );
	NAND2X1 NAND2X1_21 ( .A(target[3]), .B(H_19_), .Y(_99_) );
	OR2X2 OR2X2_4 ( .A(target[3]), .B(H_19_), .Y(_100_) );
	INVX1 INVX1_32 ( .A(target[2]), .Y(_101_) );
	NAND2X1 NAND2X1_22 ( .A(_101_), .B(_26_), .Y(_102_) );
	AOI22X1 AOI22X1_6 ( .A(_99_), .B(_100_), .C(_102_), .D(_19_), .Y(_103_) );
	INVX1 INVX1_33 ( .A(target[3]), .Y(_104_) );
	NAND2X1 NAND2X1_23 ( .A(H_19_), .B(_104_), .Y(_105_) );
	NOR2X1 NOR2X1_17 ( .A(H_19_), .B(_104_), .Y(_106_) );
	NAND2X1 NAND2X1_24 ( .A(H_18_), .B(_101_), .Y(_107_) );
	OAI21X1 OAI21X1_9 ( .A(_106_), .B(_107_), .C(_105_), .Y(_108_) );
	AOI21X1 AOI21X1_9 ( .A(_103_), .B(_98_), .C(_108_), .Y(_109_) );
	NAND2X1 NAND2X1_25 ( .A(_45_), .B(_46_), .Y(_110_) );
	NAND2X1 NAND2X1_26 ( .A(_78_), .B(_47_), .Y(_111_) );
	AOI22X1 AOI22X1_7 ( .A(_110_), .B(_30_), .C(_33_), .D(_111_), .Y(_112_) );
	NAND3X1 NAND3X1_5 ( .A(_39_), .B(_42_), .C(_112_), .Y(_113_) );
	NAND2X1 NAND2X1_27 ( .A(target[7]), .B(_46_), .Y(_114_) );
	AOI21X1 AOI21X1_10 ( .A(target[5]), .B(_40_), .C(_39_), .Y(_115_) );
	AOI22X1 AOI22X1_8 ( .A(_114_), .B(_48_), .C(_115_), .D(_112_), .Y(_116_) );
	OAI21X1 OAI21X1_10 ( .A(_109_), .B(_113_), .C(_116_), .Y(_117_) );
	NAND2X1 NAND2X1_28 ( .A(H_9_), .B(_94_), .Y(_118_) );
	OAI22X1 OAI22X1_9 ( .A(_94_), .B(H_9_), .C(H_8_), .D(_96_), .Y(_119_) );
	NAND2X1 NAND2X1_29 ( .A(_118_), .B(_119_), .Y(_120_) );
	OR2X2 OR2X2_5 ( .A(target[3]), .B(H_11_), .Y(_121_) );
	NAND2X1 NAND2X1_30 ( .A(_101_), .B(_70_), .Y(_122_) );
	AOI22X1 AOI22X1_9 ( .A(_60_), .B(_121_), .C(_122_), .D(_63_), .Y(_123_) );
	NAND2X1 NAND2X1_31 ( .A(H_11_), .B(_104_), .Y(_124_) );
	NOR2X1 NOR2X1_18 ( .A(H_11_), .B(_104_), .Y(_125_) );
	NAND2X1 NAND2X1_32 ( .A(H_10_), .B(_101_), .Y(_126_) );
	OAI21X1 OAI21X1_11 ( .A(_125_), .B(_126_), .C(_124_), .Y(_127_) );
	AOI21X1 AOI21X1_11 ( .A(_123_), .B(_120_), .C(_127_), .Y(_128_) );
	NAND2X1 NAND2X1_33 ( .A(target[6]), .B(H_14_), .Y(_129_) );
	NAND2X1 NAND2X1_34 ( .A(_78_), .B(_74_), .Y(_130_) );
	NAND2X1 NAND2X1_35 ( .A(target[7]), .B(H_15_), .Y(_131_) );
	NAND2X1 NAND2X1_36 ( .A(_45_), .B(_76_), .Y(_132_) );
	AOI22X1 AOI22X1_10 ( .A(_130_), .B(_129_), .C(_131_), .D(_132_), .Y(_133_) );
	OAI22X1 OAI22X1_10 ( .A(_37_), .B(H_13_), .C(_38_), .D(H_12_), .Y(_134_) );
	NOR2X1 NOR2X1_19 ( .A(_87_), .B(_134_), .Y(_135_) );
	NAND2X1 NAND2X1_37 ( .A(_133_), .B(_135_), .Y(_136_) );
	AOI21X1 AOI21X1_12 ( .A(target[5]), .B(_82_), .C(_81_), .Y(_137_) );
	INVX1 INVX1_34 ( .A(_1__bF_buf3), .Y(_138_) );
	NOR2X1 NOR2X1_20 ( .A(H_15_), .B(_45_), .Y(_139_) );
	OAI21X1 OAI21X1_12 ( .A(_79_), .B(_139_), .C(_138_), .Y(_140_) );
	AOI21X1 AOI21X1_13 ( .A(_133_), .B(_137_), .C(_140_), .Y(_141_) );
	OAI21X1 OAI21X1_13 ( .A(_128_), .B(_136_), .C(_141_), .Y(_142_) );
	OAI21X1 OAI21X1_14 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(bounty_synth_0_), .Y(_143_) );
	AOI21X1 AOI21X1_14 ( .A(_93_), .B(_143_), .C(_10__bF_buf6), .Y(_7__0_) );
	NAND3X1 NAND3X1_6 ( .A(H_1_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_144_) );
	OAI21X1 OAI21X1_15 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(bounty_synth_1_), .Y(_145_) );
	AOI21X1 AOI21X1_15 ( .A(_144_), .B(_145_), .C(_10__bF_buf5), .Y(_7__1_) );
	NAND3X1 NAND3X1_7 ( .A(H_2_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_146_) );
	OAI21X1 OAI21X1_16 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(bounty_synth_2_), .Y(_147_) );
	AOI21X1 AOI21X1_16 ( .A(_146_), .B(_147_), .C(_10__bF_buf4), .Y(_7__2_) );
	NAND3X1 NAND3X1_8 ( .A(H_3_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_148_) );
	OAI21X1 OAI21X1_17 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(bounty_synth_3_), .Y(_149_) );
	AOI21X1 AOI21X1_17 ( .A(_148_), .B(_149_), .C(_10__bF_buf3), .Y(_7__3_) );
	NAND3X1 NAND3X1_9 ( .A(H_4_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_150_) );
	OAI21X1 OAI21X1_18 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(bounty_synth_4_), .Y(_151_) );
	AOI21X1 AOI21X1_18 ( .A(_150_), .B(_151_), .C(_10__bF_buf2), .Y(_7__4_) );
	NAND3X1 NAND3X1_10 ( .A(H_5_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_152_) );
	OAI21X1 OAI21X1_19 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(bounty_synth_5_), .Y(_153_) );
	AOI21X1 AOI21X1_19 ( .A(_152_), .B(_153_), .C(_10__bF_buf1), .Y(_7__5_) );
	NAND3X1 NAND3X1_11 ( .A(H_6_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_154_) );
	OAI21X1 OAI21X1_20 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(bounty_synth_6_), .Y(_155_) );
	AOI21X1 AOI21X1_20 ( .A(_154_), .B(_155_), .C(_10__bF_buf0), .Y(_7__6_) );
	NAND3X1 NAND3X1_12 ( .A(H_7_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_156_) );
	OAI21X1 OAI21X1_21 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(bounty_synth_7_), .Y(_157_) );
	AOI21X1 AOI21X1_21 ( .A(_156_), .B(_157_), .C(_10__bF_buf6), .Y(_7__7_) );
	NAND3X1 NAND3X1_13 ( .A(H_8_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_158_) );
	OAI21X1 OAI21X1_22 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(bounty_synth_8_), .Y(_159_) );
	AOI21X1 AOI21X1_22 ( .A(_158_), .B(_159_), .C(_10__bF_buf5), .Y(_7__8_) );
	NAND3X1 NAND3X1_14 ( .A(H_9_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_160_) );
	OAI21X1 OAI21X1_23 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(bounty_synth_9_), .Y(_161_) );
	AOI21X1 AOI21X1_23 ( .A(_160_), .B(_161_), .C(_10__bF_buf4), .Y(_7__9_) );
	NAND3X1 NAND3X1_15 ( .A(H_10_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_162_) );
	OAI21X1 OAI21X1_24 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(bounty_synth_10_), .Y(_163_) );
	AOI21X1 AOI21X1_24 ( .A(_162_), .B(_163_), .C(_10__bF_buf3), .Y(_7__10_) );
	NAND3X1 NAND3X1_16 ( .A(H_11_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_164_) );
	OAI21X1 OAI21X1_25 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(bounty_synth_11_), .Y(_165_) );
	AOI21X1 AOI21X1_25 ( .A(_164_), .B(_165_), .C(_10__bF_buf2), .Y(_7__11_) );
	NAND3X1 NAND3X1_17 ( .A(H_12_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_166_) );
	OAI21X1 OAI21X1_26 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(bounty_synth_12_), .Y(_167_) );
	AOI21X1 AOI21X1_26 ( .A(_166_), .B(_167_), .C(_10__bF_buf1), .Y(_7__12_) );
	NAND3X1 NAND3X1_18 ( .A(H_13_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_168_) );
	OAI21X1 OAI21X1_27 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(bounty_synth_13_), .Y(_169_) );
	AOI21X1 AOI21X1_27 ( .A(_168_), .B(_169_), .C(_10__bF_buf0), .Y(_7__13_) );
	NAND3X1 NAND3X1_19 ( .A(H_14_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_170_) );
	OAI21X1 OAI21X1_28 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(bounty_synth_14_), .Y(_171_) );
	AOI21X1 AOI21X1_28 ( .A(_170_), .B(_171_), .C(_10__bF_buf6), .Y(_7__14_) );
	NAND3X1 NAND3X1_20 ( .A(H_15_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_172_) );
	OAI21X1 OAI21X1_29 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(bounty_synth_15_), .Y(_173_) );
	AOI21X1 AOI21X1_29 ( .A(_172_), .B(_173_), .C(_10__bF_buf5), .Y(_7__15_) );
	NAND3X1 NAND3X1_21 ( .A(H_16_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_174_) );
	OAI21X1 OAI21X1_30 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(bounty_synth_16_), .Y(_175_) );
	AOI21X1 AOI21X1_30 ( .A(_174_), .B(_175_), .C(_10__bF_buf4), .Y(_7__16_) );
	NAND3X1 NAND3X1_22 ( .A(H_17_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_176_) );
	OAI21X1 OAI21X1_31 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(bounty_synth_17_), .Y(_177_) );
	AOI21X1 AOI21X1_31 ( .A(_176_), .B(_177_), .C(_10__bF_buf3), .Y(_7__17_) );
	NAND3X1 NAND3X1_23 ( .A(H_18_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_178_) );
	OAI21X1 OAI21X1_32 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(bounty_synth_18_), .Y(_179_) );
	AOI21X1 AOI21X1_32 ( .A(_178_), .B(_179_), .C(_10__bF_buf2), .Y(_7__18_) );
	NAND3X1 NAND3X1_24 ( .A(H_19_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_180_) );
	OAI21X1 OAI21X1_33 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(bounty_synth_19_), .Y(_181_) );
	AOI21X1 AOI21X1_33 ( .A(_180_), .B(_181_), .C(_10__bF_buf1), .Y(_7__19_) );
	NAND3X1 NAND3X1_25 ( .A(H_20_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_182_) );
	OAI21X1 OAI21X1_34 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(bounty_synth_20_), .Y(_183_) );
	AOI21X1 AOI21X1_34 ( .A(_182_), .B(_183_), .C(_10__bF_buf0), .Y(_7__20_) );
	NAND3X1 NAND3X1_26 ( .A(H_21_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_184_) );
	OAI21X1 OAI21X1_35 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(bounty_synth_21_), .Y(_185_) );
	AOI21X1 AOI21X1_35 ( .A(_184_), .B(_185_), .C(_10__bF_buf6), .Y(_7__21_) );
	NAND3X1 NAND3X1_27 ( .A(H_22_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_186_) );
	OAI21X1 OAI21X1_36 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(bounty_synth_22_), .Y(_187_) );
	AOI21X1 AOI21X1_36 ( .A(_186_), .B(_187_), .C(_10__bF_buf5), .Y(_7__22_) );
	NAND3X1 NAND3X1_28 ( .A(H_23_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_188_) );
	OAI21X1 OAI21X1_37 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(bounty_synth_23_), .Y(_189_) );
	AOI21X1 AOI21X1_37 ( .A(_188_), .B(_189_), .C(_10__bF_buf4), .Y(_7__23_) );
	NAND3X1 NAND3X1_29 ( .A(comparador_nonce_synth_1_0_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_190_) );
	OAI21X1 OAI21X1_38 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_0_), .Y(_191_) );
	AOI21X1 AOI21X1_38 ( .A(_190_), .B(_191_), .C(_10__bF_buf3), .Y(_8__0_) );
	NAND3X1 NAND3X1_30 ( .A(comparador_nonce_synth_1_1_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_192_) );
	OAI21X1 OAI21X1_39 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_1_), .Y(_193_) );
	AOI21X1 AOI21X1_39 ( .A(_192_), .B(_193_), .C(_10__bF_buf2), .Y(_8__1_) );
	NAND3X1 NAND3X1_31 ( .A(comparador_nonce_synth_1_2_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_194_) );
	OAI21X1 OAI21X1_40 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_2_), .Y(_195_) );
	AOI21X1 AOI21X1_40 ( .A(_194_), .B(_195_), .C(_10__bF_buf1), .Y(_8__2_) );
	NAND3X1 NAND3X1_32 ( .A(comparador_nonce_synth_1_3_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_196_) );
	OAI21X1 OAI21X1_41 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_3_), .Y(_197_) );
	AOI21X1 AOI21X1_41 ( .A(_196_), .B(_197_), .C(_10__bF_buf0), .Y(_8__3_) );
	NAND3X1 NAND3X1_33 ( .A(comparador_nonce_synth_1_4_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_198_) );
	OAI21X1 OAI21X1_42 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(comparador_nonce_synth_valido_4_), .Y(_199_) );
	AOI21X1 AOI21X1_42 ( .A(_198_), .B(_199_), .C(_10__bF_buf6), .Y(_8__4_) );
	NAND3X1 NAND3X1_34 ( .A(comparador_nonce_synth_1_5_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_200_) );
	OAI21X1 OAI21X1_43 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(comparador_nonce_synth_valido_5_), .Y(_201_) );
	AOI21X1 AOI21X1_43 ( .A(_200_), .B(_201_), .C(_10__bF_buf5), .Y(_8__5_) );
	NAND3X1 NAND3X1_35 ( .A(comparador_nonce_synth_1_6_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_202_) );
	OAI21X1 OAI21X1_44 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(comparador_nonce_synth_valido_6_), .Y(_203_) );
	AOI21X1 AOI21X1_44 ( .A(_202_), .B(_203_), .C(_10__bF_buf4), .Y(_8__6_) );
	NAND3X1 NAND3X1_36 ( .A(comparador_nonce_synth_1_7_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_204_) );
	OAI21X1 OAI21X1_45 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_7_), .Y(_205_) );
	AOI21X1 AOI21X1_45 ( .A(_204_), .B(_205_), .C(_10__bF_buf3), .Y(_8__7_) );
	NAND3X1 NAND3X1_37 ( .A(comparador_nonce_synth_1_8_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_206_) );
	OAI21X1 OAI21X1_46 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_8_), .Y(_207_) );
	AOI21X1 AOI21X1_46 ( .A(_206_), .B(_207_), .C(_10__bF_buf2), .Y(_8__8_) );
	NAND3X1 NAND3X1_38 ( .A(comparador_nonce_synth_1_9_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_208_) );
	OAI21X1 OAI21X1_47 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_9_), .Y(_209_) );
	AOI21X1 AOI21X1_47 ( .A(_208_), .B(_209_), .C(_10__bF_buf1), .Y(_8__9_) );
	NAND3X1 NAND3X1_39 ( .A(comparador_nonce_synth_1_10_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_210_) );
	OAI21X1 OAI21X1_48 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_10_), .Y(_211_) );
	AOI21X1 AOI21X1_48 ( .A(_210_), .B(_211_), .C(_10__bF_buf0), .Y(_8__10_) );
	NAND3X1 NAND3X1_40 ( .A(comparador_nonce_synth_1_11_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_212_) );
	OAI21X1 OAI21X1_49 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(comparador_nonce_synth_valido_11_), .Y(_213_) );
	AOI21X1 AOI21X1_49 ( .A(_212_), .B(_213_), .C(_10__bF_buf6), .Y(_8__11_) );
	NAND3X1 NAND3X1_41 ( .A(comparador_nonce_synth_1_12_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_214_) );
	OAI21X1 OAI21X1_50 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(comparador_nonce_synth_valido_12_), .Y(_215_) );
	AOI21X1 AOI21X1_50 ( .A(_214_), .B(_215_), .C(_10__bF_buf5), .Y(_8__12_) );
	NAND3X1 NAND3X1_42 ( .A(comparador_nonce_synth_1_13_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_216_) );
	OAI21X1 OAI21X1_51 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(comparador_nonce_synth_valido_13_), .Y(_217_) );
	AOI21X1 AOI21X1_51 ( .A(_216_), .B(_217_), .C(_10__bF_buf4), .Y(_8__13_) );
	NAND3X1 NAND3X1_43 ( .A(comparador_nonce_synth_1_14_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_218_) );
	OAI21X1 OAI21X1_52 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_14_), .Y(_219_) );
	AOI21X1 AOI21X1_52 ( .A(_218_), .B(_219_), .C(_10__bF_buf3), .Y(_8__14_) );
	NAND3X1 NAND3X1_44 ( .A(comparador_nonce_synth_1_15_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_220_) );
	OAI21X1 OAI21X1_53 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_15_), .Y(_221_) );
	AOI21X1 AOI21X1_53 ( .A(_220_), .B(_221_), .C(_10__bF_buf2), .Y(_8__15_) );
	NAND3X1 NAND3X1_45 ( .A(comparador_nonce_synth_1_16_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_222_) );
	OAI21X1 OAI21X1_54 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_16_), .Y(_223_) );
	AOI21X1 AOI21X1_54 ( .A(_222_), .B(_223_), .C(_10__bF_buf1), .Y(_8__16_) );
	NAND3X1 NAND3X1_46 ( .A(comparador_nonce_synth_1_17_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_224_) );
	OAI21X1 OAI21X1_55 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_17_), .Y(_225_) );
	AOI21X1 AOI21X1_55 ( .A(_224_), .B(_225_), .C(_10__bF_buf0), .Y(_8__17_) );
	NAND3X1 NAND3X1_47 ( .A(comparador_nonce_synth_1_18_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_226_) );
	OAI21X1 OAI21X1_56 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(comparador_nonce_synth_valido_18_), .Y(_227_) );
	AOI21X1 AOI21X1_56 ( .A(_226_), .B(_227_), .C(_10__bF_buf6), .Y(_8__18_) );
	NAND3X1 NAND3X1_48 ( .A(comparador_nonce_synth_1_19_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_228_) );
	OAI21X1 OAI21X1_57 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(comparador_nonce_synth_valido_19_), .Y(_229_) );
	AOI21X1 AOI21X1_57 ( .A(_228_), .B(_229_), .C(_10__bF_buf5), .Y(_8__19_) );
	NAND3X1 NAND3X1_49 ( .A(comparador_nonce_synth_1_20_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_230_) );
	OAI21X1 OAI21X1_58 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(comparador_nonce_synth_valido_20_), .Y(_231_) );
	AOI21X1 AOI21X1_58 ( .A(_230_), .B(_231_), .C(_10__bF_buf4), .Y(_8__20_) );
	NAND3X1 NAND3X1_50 ( .A(comparador_nonce_synth_1_21_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_232_) );
	OAI21X1 OAI21X1_59 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_21_), .Y(_233_) );
	AOI21X1 AOI21X1_59 ( .A(_232_), .B(_233_), .C(_10__bF_buf3), .Y(_8__21_) );
	NAND3X1 NAND3X1_51 ( .A(comparador_nonce_synth_1_22_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_234_) );
	OAI21X1 OAI21X1_60 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_22_), .Y(_235_) );
	AOI21X1 AOI21X1_60 ( .A(_234_), .B(_235_), .C(_10__bF_buf2), .Y(_8__22_) );
	NAND3X1 NAND3X1_52 ( .A(comparador_nonce_synth_1_23_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_236_) );
	OAI21X1 OAI21X1_61 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_23_), .Y(_237_) );
	AOI21X1 AOI21X1_61 ( .A(_236_), .B(_237_), .C(_10__bF_buf1), .Y(_8__23_) );
	NAND3X1 NAND3X1_53 ( .A(comparador_nonce_synth_1_24_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_238_) );
	OAI21X1 OAI21X1_62 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_24_), .Y(_239_) );
	AOI21X1 AOI21X1_62 ( .A(_238_), .B(_239_), .C(_10__bF_buf0), .Y(_8__24_) );
	NAND3X1 NAND3X1_54 ( .A(comparador_nonce_synth_1_25_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_240_) );
	OAI21X1 OAI21X1_63 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(comparador_nonce_synth_valido_25_), .Y(_241_) );
	AOI21X1 AOI21X1_63 ( .A(_240_), .B(_241_), .C(_10__bF_buf6), .Y(_8__25_) );
	NAND3X1 NAND3X1_55 ( .A(comparador_nonce_synth_1_26_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_242_) );
	OAI21X1 OAI21X1_64 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(comparador_nonce_synth_valido_26_), .Y(_243_) );
	AOI21X1 AOI21X1_64 ( .A(_242_), .B(_243_), .C(_10__bF_buf5), .Y(_8__26_) );
	NAND3X1 NAND3X1_56 ( .A(comparador_nonce_synth_1_27_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_244_) );
	OAI21X1 OAI21X1_65 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(comparador_nonce_synth_valido_27_), .Y(_245_) );
	AOI21X1 AOI21X1_65 ( .A(_244_), .B(_245_), .C(_10__bF_buf4), .Y(_8__27_) );
	NAND3X1 NAND3X1_57 ( .A(comparador_nonce_synth_1_28_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_246_) );
	OAI21X1 OAI21X1_66 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_28_), .Y(_247_) );
	AOI21X1 AOI21X1_66 ( .A(_246_), .B(_247_), .C(_10__bF_buf3), .Y(_8__28_) );
	NAND3X1 NAND3X1_58 ( .A(comparador_nonce_synth_1_29_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_248_) );
	OAI21X1 OAI21X1_67 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_29_), .Y(_249_) );
	AOI21X1 AOI21X1_67 ( .A(_248_), .B(_249_), .C(_10__bF_buf2), .Y(_8__29_) );
	NAND3X1 NAND3X1_59 ( .A(comparador_nonce_synth_1_30_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_250_) );
	OAI21X1 OAI21X1_68 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_30_), .Y(_251_) );
	AOI21X1 AOI21X1_68 ( .A(_250_), .B(_251_), .C(_10__bF_buf1), .Y(_8__30_) );
	NAND3X1 NAND3X1_60 ( .A(comparador_nonce_synth_1_31_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_252_) );
	OAI21X1 OAI21X1_69 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_31_), .Y(_253_) );
	AOI21X1 AOI21X1_69 ( .A(_252_), .B(_253_), .C(_10__bF_buf0), .Y(_8__31_) );
	AOI21X1 AOI21X1_70 ( .A(_53__bF_buf6), .B(_92__bF_buf6), .C(comparador_valid_bF_buf5), .Y(_254_) );
	OAI21X1 OAI21X1_70 ( .A(_53__bF_buf5), .B(_1__bF_buf2), .C(reset_L_bF_buf5), .Y(_255_) );
	NOR2X1 NOR2X1_21 ( .A(_255_), .B(_254_), .Y(_9_) );
	DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf62), .D(_9_), .Q(comparador_valid) );
	DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf61), .D(_8__0_), .Q(comparador_nonce_synth_valido_0_) );
	DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf60), .D(_8__1_), .Q(comparador_nonce_synth_valido_1_) );
	DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf59), .D(_8__2_), .Q(comparador_nonce_synth_valido_2_) );
	DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf58), .D(_8__3_), .Q(comparador_nonce_synth_valido_3_) );
	DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf57), .D(_8__4_), .Q(comparador_nonce_synth_valido_4_) );
	DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf56), .D(_8__5_), .Q(comparador_nonce_synth_valido_5_) );
	DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf55), .D(_8__6_), .Q(comparador_nonce_synth_valido_6_) );
	DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf54), .D(_8__7_), .Q(comparador_nonce_synth_valido_7_) );
	DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf53), .D(_8__8_), .Q(comparador_nonce_synth_valido_8_) );
	DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf52), .D(_8__9_), .Q(comparador_nonce_synth_valido_9_) );
	DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf51), .D(_8__10_), .Q(comparador_nonce_synth_valido_10_) );
	DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf50), .D(_8__11_), .Q(comparador_nonce_synth_valido_11_) );
	DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf49), .D(_8__12_), .Q(comparador_nonce_synth_valido_12_) );
	DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf48), .D(_8__13_), .Q(comparador_nonce_synth_valido_13_) );
	DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf47), .D(_8__14_), .Q(comparador_nonce_synth_valido_14_) );
	DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf46), .D(_8__15_), .Q(comparador_nonce_synth_valido_15_) );
	DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf45), .D(_8__16_), .Q(comparador_nonce_synth_valido_16_) );
	DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf44), .D(_8__17_), .Q(comparador_nonce_synth_valido_17_) );
	DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf43), .D(_8__18_), .Q(comparador_nonce_synth_valido_18_) );
	DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf42), .D(_8__19_), .Q(comparador_nonce_synth_valido_19_) );
	DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf41), .D(_8__20_), .Q(comparador_nonce_synth_valido_20_) );
	DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf40), .D(_8__21_), .Q(comparador_nonce_synth_valido_21_) );
	DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf39), .D(_8__22_), .Q(comparador_nonce_synth_valido_22_) );
	DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf38), .D(_8__23_), .Q(comparador_nonce_synth_valido_23_) );
	DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf37), .D(_8__24_), .Q(comparador_nonce_synth_valido_24_) );
	DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf36), .D(_8__25_), .Q(comparador_nonce_synth_valido_25_) );
	DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf35), .D(_8__26_), .Q(comparador_nonce_synth_valido_26_) );
	DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf34), .D(_8__27_), .Q(comparador_nonce_synth_valido_27_) );
	DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf33), .D(_8__28_), .Q(comparador_nonce_synth_valido_28_) );
	DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf32), .D(_8__29_), .Q(comparador_nonce_synth_valido_29_) );
	DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf31), .D(_8__30_), .Q(comparador_nonce_synth_valido_30_) );
	DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf30), .D(_8__31_), .Q(comparador_nonce_synth_valido_31_) );
	DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf29), .D(_7__0_), .Q(bounty_synth_0_) );
	DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf28), .D(_7__1_), .Q(bounty_synth_1_) );
	DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf27), .D(_7__2_), .Q(bounty_synth_2_) );
	DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf26), .D(_7__3_), .Q(bounty_synth_3_) );
	DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf25), .D(_7__4_), .Q(bounty_synth_4_) );
	DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf24), .D(_7__5_), .Q(bounty_synth_5_) );
	DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf23), .D(_7__6_), .Q(bounty_synth_6_) );
	DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf22), .D(_7__7_), .Q(bounty_synth_7_) );
	DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf21), .D(_7__8_), .Q(bounty_synth_8_) );
	DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf20), .D(_7__9_), .Q(bounty_synth_9_) );
	DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf19), .D(_7__10_), .Q(bounty_synth_10_) );
	DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf18), .D(_7__11_), .Q(bounty_synth_11_) );
	DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf17), .D(_7__12_), .Q(bounty_synth_12_) );
	DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf16), .D(_7__13_), .Q(bounty_synth_13_) );
	DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf15), .D(_7__14_), .Q(bounty_synth_14_) );
	DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf14), .D(_7__15_), .Q(bounty_synth_15_) );
	DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf13), .D(_7__16_), .Q(bounty_synth_16_) );
	DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf12), .D(_7__17_), .Q(bounty_synth_17_) );
	DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf11), .D(_7__18_), .Q(bounty_synth_18_) );
	DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf10), .D(_7__19_), .Q(bounty_synth_19_) );
	DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf9), .D(_7__20_), .Q(bounty_synth_20_) );
	DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf8), .D(_7__21_), .Q(bounty_synth_21_) );
	DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf7), .D(_7__22_), .Q(bounty_synth_22_) );
	DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf6), .D(_7__23_), .Q(bounty_synth_23_) );
	INVX1 INVX1_35 ( .A(bloque_in_32_), .Y(_257_) );
	NOR2X1 NOR2X1_22 ( .A(concatenador_count_1_bF_buf6), .B(concatenador_count_0_bF_buf11), .Y(_258_) );
	NOR2X1 NOR2X1_23 ( .A(concatenador_count_3_), .B(concatenador_count_2_), .Y(_259_) );
	NOR2X1 NOR2X1_24 ( .A(concatenador_count_5_), .B(concatenador_count_4_), .Y(_260_) );
	NAND3X1 NAND3X1_61 ( .A(_258_), .B(_259_), .C(_260_), .Y(_261_) );
	OAI21X1 OAI21X1_71 ( .A(_261__bF_buf15), .B(RAM_entrada_89_), .C(reset_L_bF_buf4), .Y(_262_) );
	AOI21X1 AOI21X1_71 ( .A(_257_), .B(_261__bF_buf14), .C(_262_), .Y(_256__32_) );
	INVX1 INVX1_36 ( .A(bloque_in_33_), .Y(_263_) );
	OAI21X1 OAI21X1_72 ( .A(_261__bF_buf13), .B(RAM_entrada_77_), .C(reset_L_bF_buf3), .Y(_264_) );
	AOI21X1 AOI21X1_72 ( .A(_263_), .B(_261__bF_buf12), .C(_264_), .Y(_256__33_) );
	INVX1 INVX1_37 ( .A(bloque_in_34_), .Y(_265_) );
	OAI21X1 OAI21X1_73 ( .A(_261__bF_buf11), .B(RAM_entrada_84_), .C(reset_L_bF_buf2), .Y(_266_) );
	AOI21X1 AOI21X1_73 ( .A(_265_), .B(_261__bF_buf10), .C(_266_), .Y(_256__34_) );
	INVX1 INVX1_38 ( .A(bloque_in_35_), .Y(_267_) );
	OAI21X1 OAI21X1_74 ( .A(_261__bF_buf9), .B(RAM_entrada_94_), .C(reset_L_bF_buf1), .Y(_268_) );
	AOI21X1 AOI21X1_74 ( .A(_267_), .B(_261__bF_buf8), .C(_268_), .Y(_256__35_) );
	INVX1 INVX1_39 ( .A(bloque_in_36_), .Y(_269_) );
	OAI21X1 OAI21X1_75 ( .A(_261__bF_buf7), .B(RAM_entrada_94_), .C(reset_L_bF_buf0), .Y(_270_) );
	AOI21X1 AOI21X1_75 ( .A(_269_), .B(_261__bF_buf6), .C(_270_), .Y(_256__36_) );
	INVX1 INVX1_40 ( .A(bloque_in_37_), .Y(_271_) );
	OAI21X1 OAI21X1_76 ( .A(_261__bF_buf5), .B(RAM_entrada_93_), .C(reset_L_bF_buf11), .Y(_272_) );
	AOI21X1 AOI21X1_76 ( .A(_271_), .B(_261__bF_buf4), .C(_272_), .Y(_256__37_) );
	INVX1 INVX1_41 ( .A(bloque_in_38_), .Y(_273_) );
	OAI21X1 OAI21X1_77 ( .A(_261__bF_buf3), .B(RAM_entrada_95_), .C(reset_L_bF_buf10), .Y(_274_) );
	AOI21X1 AOI21X1_77 ( .A(_273_), .B(_261__bF_buf2), .C(_274_), .Y(_256__38_) );
	INVX1 INVX1_42 ( .A(bloque_in_39_), .Y(_275_) );
	OAI21X1 OAI21X1_78 ( .A(_261__bF_buf1), .B(RAM_entrada_95_), .C(reset_L_bF_buf9), .Y(_276_) );
	AOI21X1 AOI21X1_78 ( .A(_275_), .B(_261__bF_buf0), .C(_276_), .Y(_256__39_) );
	INVX1 INVX1_43 ( .A(bloque_in_40_), .Y(_277_) );
	OAI21X1 OAI21X1_79 ( .A(_261__bF_buf15), .B(RAM_entrada_86_), .C(reset_L_bF_buf8), .Y(_278_) );
	AOI21X1 AOI21X1_79 ( .A(_277_), .B(_261__bF_buf14), .C(_278_), .Y(_256__40_) );
	INVX1 INVX1_44 ( .A(bloque_in_41_), .Y(_279_) );
	OAI21X1 OAI21X1_80 ( .A(_261__bF_buf13), .B(RAM_entrada_84_), .C(reset_L_bF_buf7), .Y(_280_) );
	AOI21X1 AOI21X1_80 ( .A(_279_), .B(_261__bF_buf12), .C(_280_), .Y(_256__41_) );
	INVX1 INVX1_45 ( .A(bloque_in_42_), .Y(_281_) );
	OAI21X1 OAI21X1_81 ( .A(_261__bF_buf11), .B(RAM_entrada_77_), .C(reset_L_bF_buf6), .Y(_282_) );
	AOI21X1 AOI21X1_81 ( .A(_281_), .B(_261__bF_buf10), .C(_282_), .Y(_256__42_) );
	INVX1 INVX1_46 ( .A(bloque_in_43_), .Y(_283_) );
	OAI21X1 OAI21X1_82 ( .A(_261__bF_buf9), .B(RAM_entrada_46_), .C(reset_L_bF_buf5), .Y(_284_) );
	AOI21X1 AOI21X1_82 ( .A(_283_), .B(_261__bF_buf8), .C(_284_), .Y(_256__43_) );
	INVX1 INVX1_47 ( .A(bloque_in_44_), .Y(_285_) );
	OAI21X1 OAI21X1_83 ( .A(_261__bF_buf7), .B(RAM_entrada_82_), .C(reset_L_bF_buf4), .Y(_286_) );
	AOI21X1 AOI21X1_83 ( .A(_285_), .B(_261__bF_buf6), .C(_286_), .Y(_256__44_) );
	INVX1 INVX1_48 ( .A(bloque_in_45_), .Y(_287_) );
	OAI21X1 OAI21X1_84 ( .A(_261__bF_buf5), .B(RAM_entrada_92_), .C(reset_L_bF_buf3), .Y(_288_) );
	AOI21X1 AOI21X1_84 ( .A(_287_), .B(_261__bF_buf4), .C(_288_), .Y(_256__45_) );
	INVX1 INVX1_49 ( .A(bloque_in_46_), .Y(_289_) );
	OAI21X1 OAI21X1_85 ( .A(_261__bF_buf3), .B(RAM_entrada_71_), .C(reset_L_bF_buf2), .Y(_290_) );
	AOI21X1 AOI21X1_85 ( .A(_289_), .B(_261__bF_buf2), .C(_290_), .Y(_256__46_) );
	INVX1 INVX1_50 ( .A(bloque_in_47_), .Y(_291_) );
	OAI21X1 OAI21X1_86 ( .A(_261__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf1), .Y(_292_) );
	AOI21X1 AOI21X1_86 ( .A(_291_), .B(_261__bF_buf0), .C(_292_), .Y(_256__47_) );
	INVX1 INVX1_51 ( .A(bloque_in_48_), .Y(_293_) );
	OAI21X1 OAI21X1_87 ( .A(_261__bF_buf15), .B(RAM_entrada_92_), .C(reset_L_bF_buf0), .Y(_294_) );
	AOI21X1 AOI21X1_87 ( .A(_293_), .B(_261__bF_buf14), .C(_294_), .Y(_256__48_) );
	INVX1 INVX1_52 ( .A(bloque_in_49_), .Y(_295_) );
	OAI21X1 OAI21X1_88 ( .A(_261__bF_buf13), .B(RAM_entrada_84_), .C(reset_L_bF_buf11), .Y(_296_) );
	AOI21X1 AOI21X1_88 ( .A(_295_), .B(_261__bF_buf12), .C(_296_), .Y(_256__49_) );
	INVX1 INVX1_53 ( .A(bloque_in_50_), .Y(_297_) );
	OAI21X1 OAI21X1_89 ( .A(_261__bF_buf11), .B(RAM_entrada_86_), .C(reset_L_bF_buf10), .Y(_298_) );
	AOI21X1 AOI21X1_89 ( .A(_297_), .B(_261__bF_buf10), .C(_298_), .Y(_256__50_) );
	INVX1 INVX1_54 ( .A(bloque_in_51_), .Y(_299_) );
	OAI21X1 OAI21X1_90 ( .A(_261__bF_buf9), .B(RAM_entrada_86_), .C(reset_L_bF_buf9), .Y(_300_) );
	AOI21X1 AOI21X1_90 ( .A(_299_), .B(_261__bF_buf8), .C(_300_), .Y(_256__51_) );
	INVX1 INVX1_55 ( .A(bloque_in_52_), .Y(_301_) );
	OAI21X1 OAI21X1_91 ( .A(_261__bF_buf7), .B(vdd), .C(reset_L_bF_buf8), .Y(_302_) );
	AOI21X1 AOI21X1_91 ( .A(_301_), .B(_261__bF_buf6), .C(_302_), .Y(_256__52_) );
	INVX1 INVX1_56 ( .A(bloque_in_53_), .Y(_303_) );
	OAI21X1 OAI21X1_92 ( .A(_261__bF_buf5), .B(RAM_entrada_58_), .C(reset_L_bF_buf7), .Y(_304_) );
	AOI21X1 AOI21X1_92 ( .A(_303_), .B(_261__bF_buf4), .C(_304_), .Y(_256__53_) );
	INVX1 INVX1_57 ( .A(bloque_in_54_), .Y(_305_) );
	OAI21X1 OAI21X1_93 ( .A(_261__bF_buf3), .B(gnd), .C(reset_L_bF_buf6), .Y(_306_) );
	AOI21X1 AOI21X1_93 ( .A(_305_), .B(_261__bF_buf2), .C(_306_), .Y(_256__54_) );
	INVX1 INVX1_58 ( .A(bloque_in_55_), .Y(_307_) );
	OAI21X1 OAI21X1_94 ( .A(_261__bF_buf1), .B(RAM_entrada_71_), .C(reset_L_bF_buf5), .Y(_308_) );
	AOI21X1 AOI21X1_94 ( .A(_307_), .B(_261__bF_buf0), .C(_308_), .Y(_256__55_) );
	INVX1 INVX1_59 ( .A(bloque_in_56_), .Y(_309_) );
	OAI21X1 OAI21X1_95 ( .A(_261__bF_buf15), .B(RAM_entrada_88_), .C(reset_L_bF_buf4), .Y(_310_) );
	AOI21X1 AOI21X1_95 ( .A(_309_), .B(_261__bF_buf14), .C(_310_), .Y(_256__56_) );
	INVX1 INVX1_60 ( .A(bloque_in_57_), .Y(_311_) );
	OAI21X1 OAI21X1_96 ( .A(_261__bF_buf13), .B(RAM_entrada_93_), .C(reset_L_bF_buf3), .Y(_312_) );
	AOI21X1 AOI21X1_96 ( .A(_311_), .B(_261__bF_buf12), .C(_312_), .Y(_256__57_) );
	INVX1 INVX1_61 ( .A(bloque_in_58_), .Y(_313_) );
	OAI21X1 OAI21X1_97 ( .A(_261__bF_buf11), .B(RAM_entrada_58_), .C(reset_L_bF_buf2), .Y(_314_) );
	AOI21X1 AOI21X1_97 ( .A(_313_), .B(_261__bF_buf10), .C(_314_), .Y(_256__58_) );
	INVX1 INVX1_62 ( .A(bloque_in_59_), .Y(_315_) );
	OAI21X1 OAI21X1_98 ( .A(_261__bF_buf9), .B(RAM_entrada_85_), .C(reset_L_bF_buf1), .Y(_316_) );
	AOI21X1 AOI21X1_98 ( .A(_315_), .B(_261__bF_buf8), .C(_316_), .Y(_256__59_) );
	INVX1 INVX1_63 ( .A(bloque_in_60_), .Y(_317_) );
	OAI21X1 OAI21X1_99 ( .A(_261__bF_buf7), .B(RAM_entrada_71_), .C(reset_L_bF_buf0), .Y(_318_) );
	AOI21X1 AOI21X1_99 ( .A(_317_), .B(_261__bF_buf6), .C(_318_), .Y(_256__60_) );
	INVX1 INVX1_64 ( .A(bloque_in_61_), .Y(_319_) );
	OAI21X1 OAI21X1_100 ( .A(_261__bF_buf5), .B(RAM_entrada_93_), .C(reset_L_bF_buf11), .Y(_320_) );
	AOI21X1 AOI21X1_100 ( .A(_319_), .B(_261__bF_buf4), .C(_320_), .Y(_256__61_) );
	INVX1 INVX1_65 ( .A(bloque_in_62_), .Y(_321_) );
	OAI21X1 OAI21X1_101 ( .A(_261__bF_buf3), .B(RAM_entrada_84_), .C(reset_L_bF_buf10), .Y(_322_) );
	AOI21X1 AOI21X1_101 ( .A(_321_), .B(_261__bF_buf2), .C(_322_), .Y(_256__62_) );
	INVX1 INVX1_66 ( .A(bloque_in_63_), .Y(_323_) );
	OAI21X1 OAI21X1_102 ( .A(_261__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf9), .Y(_324_) );
	AOI21X1 AOI21X1_102 ( .A(_323_), .B(_261__bF_buf0), .C(_324_), .Y(_256__63_) );
	INVX1 INVX1_67 ( .A(bloque_in_64_), .Y(_325_) );
	OAI21X1 OAI21X1_103 ( .A(_261__bF_buf15), .B(RAM_entrada_71_), .C(reset_L_bF_buf8), .Y(_326_) );
	AOI21X1 AOI21X1_103 ( .A(_325_), .B(_261__bF_buf14), .C(_326_), .Y(_256__64_) );
	INVX1 INVX1_68 ( .A(bloque_in_65_), .Y(_327_) );
	OAI21X1 OAI21X1_104 ( .A(_261__bF_buf13), .B(RAM_entrada_95_), .C(reset_L_bF_buf7), .Y(_328_) );
	AOI21X1 AOI21X1_104 ( .A(_327_), .B(_261__bF_buf12), .C(_328_), .Y(_256__65_) );
	INVX1 INVX1_69 ( .A(bloque_in_66_), .Y(_329_) );
	OAI21X1 OAI21X1_105 ( .A(_261__bF_buf11), .B(RAM_entrada_92_), .C(reset_L_bF_buf6), .Y(_330_) );
	AOI21X1 AOI21X1_105 ( .A(_329_), .B(_261__bF_buf10), .C(_330_), .Y(_256__66_) );
	INVX1 INVX1_70 ( .A(bloque_in_67_), .Y(_331_) );
	OAI21X1 OAI21X1_106 ( .A(_261__bF_buf9), .B(RAM_entrada_92_), .C(reset_L_bF_buf5), .Y(_332_) );
	AOI21X1 AOI21X1_106 ( .A(_331_), .B(_261__bF_buf8), .C(_332_), .Y(_256__67_) );
	INVX1 INVX1_71 ( .A(bloque_in_68_), .Y(_333_) );
	OAI21X1 OAI21X1_107 ( .A(_261__bF_buf7), .B(RAM_entrada_71_), .C(reset_L_bF_buf4), .Y(_334_) );
	AOI21X1 AOI21X1_107 ( .A(_333_), .B(_261__bF_buf6), .C(_334_), .Y(_256__68_) );
	INVX1 INVX1_72 ( .A(bloque_in_69_), .Y(_335_) );
	OAI21X1 OAI21X1_108 ( .A(_261__bF_buf5), .B(RAM_entrada_84_), .C(reset_L_bF_buf3), .Y(_336_) );
	AOI21X1 AOI21X1_108 ( .A(_335_), .B(_261__bF_buf4), .C(_336_), .Y(_256__69_) );
	INVX1 INVX1_73 ( .A(bloque_in_70_), .Y(_337_) );
	OAI21X1 OAI21X1_109 ( .A(_261__bF_buf3), .B(RAM_entrada_84_), .C(reset_L_bF_buf2), .Y(_338_) );
	AOI21X1 AOI21X1_109 ( .A(_337_), .B(_261__bF_buf2), .C(_338_), .Y(_256__70_) );
	INVX1 INVX1_74 ( .A(bloque_in_71_), .Y(_339_) );
	OAI21X1 OAI21X1_110 ( .A(_261__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf1), .Y(_340_) );
	AOI21X1 AOI21X1_110 ( .A(_339_), .B(_261__bF_buf0), .C(_340_), .Y(_256__71_) );
	INVX1 INVX1_75 ( .A(bloque_in_72_), .Y(_341_) );
	OAI21X1 OAI21X1_111 ( .A(_261__bF_buf15), .B(RAM_entrada_89_), .C(reset_L_bF_buf0), .Y(_342_) );
	AOI21X1 AOI21X1_111 ( .A(_341_), .B(_261__bF_buf14), .C(_342_), .Y(_256__72_) );
	INVX1 INVX1_76 ( .A(bloque_in_73_), .Y(_343_) );
	OAI21X1 OAI21X1_112 ( .A(_261__bF_buf13), .B(RAM_entrada_82_), .C(reset_L_bF_buf11), .Y(_344_) );
	AOI21X1 AOI21X1_112 ( .A(_343_), .B(_261__bF_buf12), .C(_344_), .Y(_256__73_) );
	INVX1 INVX1_77 ( .A(bloque_in_74_), .Y(_345_) );
	OAI21X1 OAI21X1_113 ( .A(_261__bF_buf11), .B(RAM_entrada_92_), .C(reset_L_bF_buf10), .Y(_346_) );
	AOI21X1 AOI21X1_113 ( .A(_345_), .B(_261__bF_buf10), .C(_346_), .Y(_256__74_) );
	INVX1 INVX1_78 ( .A(bloque_in_75_), .Y(_347_) );
	OAI21X1 OAI21X1_114 ( .A(_261__bF_buf9), .B(RAM_entrada_85_), .C(reset_L_bF_buf9), .Y(_348_) );
	AOI21X1 AOI21X1_114 ( .A(_347_), .B(_261__bF_buf8), .C(_348_), .Y(_256__75_) );
	INVX1 INVX1_79 ( .A(bloque_in_76_), .Y(_349_) );
	OAI21X1 OAI21X1_115 ( .A(_261__bF_buf7), .B(RAM_entrada_82_), .C(reset_L_bF_buf8), .Y(_350_) );
	AOI21X1 AOI21X1_115 ( .A(_349_), .B(_261__bF_buf6), .C(_350_), .Y(_256__76_) );
	INVX1 INVX1_80 ( .A(bloque_in_77_), .Y(_351_) );
	OAI21X1 OAI21X1_116 ( .A(_261__bF_buf5), .B(RAM_entrada_46_), .C(reset_L_bF_buf7), .Y(_352_) );
	AOI21X1 AOI21X1_116 ( .A(_351_), .B(_261__bF_buf4), .C(_352_), .Y(_256__77_) );
	INVX1 INVX1_81 ( .A(bloque_in_78_), .Y(_353_) );
	OAI21X1 OAI21X1_117 ( .A(_261__bF_buf3), .B(RAM_entrada_46_), .C(reset_L_bF_buf6), .Y(_354_) );
	AOI21X1 AOI21X1_117 ( .A(_353_), .B(_261__bF_buf2), .C(_354_), .Y(_256__78_) );
	INVX1 INVX1_82 ( .A(bloque_in_79_), .Y(_355_) );
	OAI21X1 OAI21X1_118 ( .A(_261__bF_buf1), .B(vdd), .C(reset_L_bF_buf5), .Y(_356_) );
	AOI21X1 AOI21X1_118 ( .A(_355_), .B(_261__bF_buf0), .C(_356_), .Y(_256__79_) );
	INVX1 INVX1_83 ( .A(bloque_in_80_), .Y(_357_) );
	OAI21X1 OAI21X1_119 ( .A(_261__bF_buf15), .B(RAM_entrada_71_), .C(reset_L_bF_buf4), .Y(_358_) );
	AOI21X1 AOI21X1_119 ( .A(_357_), .B(_261__bF_buf14), .C(_358_), .Y(_256__80_) );
	INVX1 INVX1_84 ( .A(bloque_in_81_), .Y(_359_) );
	OAI21X1 OAI21X1_120 ( .A(_261__bF_buf13), .B(RAM_entrada_84_), .C(reset_L_bF_buf3), .Y(_360_) );
	AOI21X1 AOI21X1_120 ( .A(_359_), .B(_261__bF_buf12), .C(_360_), .Y(_256__81_) );
	INVX1 INVX1_85 ( .A(bloque_in_82_), .Y(_361_) );
	OAI21X1 OAI21X1_121 ( .A(_261__bF_buf11), .B(RAM_entrada_71_), .C(reset_L_bF_buf2), .Y(_362_) );
	AOI21X1 AOI21X1_121 ( .A(_361_), .B(_261__bF_buf10), .C(_362_), .Y(_256__82_) );
	INVX1 INVX1_86 ( .A(bloque_in_83_), .Y(_363_) );
	OAI21X1 OAI21X1_122 ( .A(_261__bF_buf9), .B(RAM_entrada_93_), .C(reset_L_bF_buf1), .Y(_364_) );
	AOI21X1 AOI21X1_122 ( .A(_363_), .B(_261__bF_buf8), .C(_364_), .Y(_256__83_) );
	INVX1 INVX1_87 ( .A(bloque_in_84_), .Y(_365_) );
	OAI21X1 OAI21X1_123 ( .A(_261__bF_buf7), .B(RAM_entrada_89_), .C(reset_L_bF_buf0), .Y(_366_) );
	AOI21X1 AOI21X1_123 ( .A(_365_), .B(_261__bF_buf6), .C(_366_), .Y(_256__84_) );
	INVX1 INVX1_88 ( .A(bloque_in_85_), .Y(_367_) );
	OAI21X1 OAI21X1_124 ( .A(_261__bF_buf5), .B(RAM_entrada_71_), .C(reset_L_bF_buf11), .Y(_368_) );
	AOI21X1 AOI21X1_124 ( .A(_367_), .B(_261__bF_buf4), .C(_368_), .Y(_256__85_) );
	INVX1 INVX1_89 ( .A(bloque_in_86_), .Y(_369_) );
	OAI21X1 OAI21X1_125 ( .A(_261__bF_buf3), .B(RAM_entrada_84_), .C(reset_L_bF_buf10), .Y(_370_) );
	AOI21X1 AOI21X1_125 ( .A(_369_), .B(_261__bF_buf2), .C(_370_), .Y(_256__86_) );
	INVX1 INVX1_90 ( .A(bloque_in_87_), .Y(_371_) );
	OAI21X1 OAI21X1_126 ( .A(_261__bF_buf1), .B(RAM_entrada_85_), .C(reset_L_bF_buf9), .Y(_372_) );
	AOI21X1 AOI21X1_126 ( .A(_371_), .B(_261__bF_buf0), .C(_372_), .Y(_256__87_) );
	INVX1 INVX1_91 ( .A(bloque_in_88_), .Y(_373_) );
	OAI21X1 OAI21X1_127 ( .A(_261__bF_buf15), .B(RAM_entrada_89_), .C(reset_L_bF_buf8), .Y(_374_) );
	AOI21X1 AOI21X1_127 ( .A(_373_), .B(_261__bF_buf14), .C(_374_), .Y(_256__88_) );
	INVX1 INVX1_92 ( .A(bloque_in_89_), .Y(_375_) );
	OAI21X1 OAI21X1_128 ( .A(_261__bF_buf13), .B(RAM_entrada_58_), .C(reset_L_bF_buf7), .Y(_376_) );
	AOI21X1 AOI21X1_128 ( .A(_375_), .B(_261__bF_buf12), .C(_376_), .Y(_256__89_) );
	INVX1 INVX1_93 ( .A(bloque_in_90_), .Y(_377_) );
	OAI21X1 OAI21X1_129 ( .A(_261__bF_buf11), .B(RAM_entrada_58_), .C(reset_L_bF_buf6), .Y(_378_) );
	AOI21X1 AOI21X1_129 ( .A(_377_), .B(_261__bF_buf10), .C(_378_), .Y(_256__90_) );
	INVX1 INVX1_94 ( .A(bloque_in_91_), .Y(_379_) );
	OAI21X1 OAI21X1_130 ( .A(_261__bF_buf9), .B(RAM_entrada_95_), .C(reset_L_bF_buf5), .Y(_380_) );
	AOI21X1 AOI21X1_130 ( .A(_379_), .B(_261__bF_buf8), .C(_380_), .Y(_256__91_) );
	INVX1 INVX1_95 ( .A(bloque_in_92_), .Y(_381_) );
	OAI21X1 OAI21X1_131 ( .A(_261__bF_buf7), .B(RAM_entrada_94_), .C(reset_L_bF_buf4), .Y(_382_) );
	AOI21X1 AOI21X1_131 ( .A(_381_), .B(_261__bF_buf6), .C(_382_), .Y(_256__92_) );
	INVX1 INVX1_96 ( .A(bloque_in_93_), .Y(_383_) );
	OAI21X1 OAI21X1_132 ( .A(_261__bF_buf5), .B(RAM_entrada_71_), .C(reset_L_bF_buf3), .Y(_384_) );
	AOI21X1 AOI21X1_132 ( .A(_383_), .B(_261__bF_buf4), .C(_384_), .Y(_256__93_) );
	INVX1 INVX1_97 ( .A(bloque_in_94_), .Y(_385_) );
	OAI21X1 OAI21X1_133 ( .A(_261__bF_buf3), .B(RAM_entrada_86_), .C(reset_L_bF_buf2), .Y(_386_) );
	AOI21X1 AOI21X1_133 ( .A(_385_), .B(_261__bF_buf2), .C(_386_), .Y(_256__94_) );
	INVX1 INVX1_98 ( .A(bloque_in_95_), .Y(_387_) );
	OAI21X1 OAI21X1_134 ( .A(_261__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf1), .Y(_388_) );
	AOI21X1 AOI21X1_134 ( .A(_387_), .B(_261__bF_buf0), .C(_388_), .Y(_256__95_) );
	INVX1 INVX1_99 ( .A(bloque_in_96_), .Y(_389_) );
	OAI21X1 OAI21X1_135 ( .A(_261__bF_buf15), .B(RAM_entrada_88_), .C(reset_L_bF_buf0), .Y(_390_) );
	AOI21X1 AOI21X1_135 ( .A(_389_), .B(_261__bF_buf14), .C(_390_), .Y(_256__96_) );
	INVX1 INVX1_100 ( .A(bloque_in_97_), .Y(_391_) );
	OAI21X1 OAI21X1_136 ( .A(_261__bF_buf13), .B(RAM_entrada_93_), .C(reset_L_bF_buf11), .Y(_392_) );
	AOI21X1 AOI21X1_136 ( .A(_391_), .B(_261__bF_buf12), .C(_392_), .Y(_256__97_) );
	INVX1 INVX1_101 ( .A(bloque_in_98_), .Y(_393_) );
	OAI21X1 OAI21X1_137 ( .A(_261__bF_buf11), .B(RAM_entrada_93_), .C(reset_L_bF_buf10), .Y(_394_) );
	AOI21X1 AOI21X1_137 ( .A(_393_), .B(_261__bF_buf10), .C(_394_), .Y(_256__98_) );
	INVX1 INVX1_102 ( .A(bloque_in_99_), .Y(_395_) );
	OAI21X1 OAI21X1_138 ( .A(_261__bF_buf9), .B(vdd), .C(reset_L_bF_buf9), .Y(_396_) );
	AOI21X1 AOI21X1_138 ( .A(_395_), .B(_261__bF_buf8), .C(_396_), .Y(_256__99_) );
	INVX1 INVX1_103 ( .A(bloque_in_100_), .Y(_397_) );
	OAI21X1 OAI21X1_139 ( .A(_261__bF_buf7), .B(RAM_entrada_89_), .C(reset_L_bF_buf8), .Y(_398_) );
	AOI21X1 AOI21X1_139 ( .A(_397_), .B(_261__bF_buf6), .C(_398_), .Y(_256__100_) );
	INVX1 INVX1_104 ( .A(bloque_in_101_), .Y(_399_) );
	OAI21X1 OAI21X1_140 ( .A(_261__bF_buf5), .B(RAM_entrada_82_), .C(reset_L_bF_buf7), .Y(_400_) );
	AOI21X1 AOI21X1_140 ( .A(_399_), .B(_261__bF_buf4), .C(_400_), .Y(_256__101_) );
	INVX1 INVX1_105 ( .A(bloque_in_102_), .Y(_401_) );
	OAI21X1 OAI21X1_141 ( .A(_261__bF_buf3), .B(RAM_entrada_71_), .C(reset_L_bF_buf6), .Y(_402_) );
	AOI21X1 AOI21X1_141 ( .A(_401_), .B(_261__bF_buf2), .C(_402_), .Y(_256__102_) );
	INVX1 INVX1_106 ( .A(bloque_in_103_), .Y(_403_) );
	OAI21X1 OAI21X1_142 ( .A(_261__bF_buf1), .B(RAM_entrada_71_), .C(reset_L_bF_buf5), .Y(_404_) );
	AOI21X1 AOI21X1_142 ( .A(_403_), .B(_261__bF_buf0), .C(_404_), .Y(_256__103_) );
	INVX1 INVX1_107 ( .A(bloque_in_104_), .Y(_405_) );
	OAI21X1 OAI21X1_143 ( .A(_261__bF_buf15), .B(RAM_entrada_92_), .C(reset_L_bF_buf4), .Y(_406_) );
	AOI21X1 AOI21X1_143 ( .A(_405_), .B(_261__bF_buf14), .C(_406_), .Y(_256__104_) );
	INVX1 INVX1_108 ( .A(bloque_in_105_), .Y(_407_) );
	OAI21X1 OAI21X1_144 ( .A(_261__bF_buf13), .B(RAM_entrada_88_), .C(reset_L_bF_buf3), .Y(_408_) );
	AOI21X1 AOI21X1_144 ( .A(_407_), .B(_261__bF_buf12), .C(_408_), .Y(_256__105_) );
	INVX1 INVX1_109 ( .A(bloque_in_106_), .Y(_409_) );
	OAI21X1 OAI21X1_145 ( .A(_261__bF_buf11), .B(RAM_entrada_88_), .C(reset_L_bF_buf2), .Y(_410_) );
	AOI21X1 AOI21X1_145 ( .A(_409_), .B(_261__bF_buf10), .C(_410_), .Y(_256__106_) );
	INVX1 INVX1_110 ( .A(bloque_in_107_), .Y(_411_) );
	OAI21X1 OAI21X1_146 ( .A(_261__bF_buf9), .B(vdd), .C(reset_L_bF_buf1), .Y(_412_) );
	AOI21X1 AOI21X1_146 ( .A(_411_), .B(_261__bF_buf8), .C(_412_), .Y(_256__107_) );
	INVX1 INVX1_111 ( .A(bloque_in_108_), .Y(_413_) );
	OAI21X1 OAI21X1_147 ( .A(_261__bF_buf7), .B(RAM_entrada_84_), .C(reset_L_bF_buf0), .Y(_414_) );
	AOI21X1 AOI21X1_147 ( .A(_413_), .B(_261__bF_buf6), .C(_414_), .Y(_256__108_) );
	INVX1 INVX1_112 ( .A(bloque_in_109_), .Y(_415_) );
	OAI21X1 OAI21X1_148 ( .A(_261__bF_buf5), .B(RAM_entrada_77_), .C(reset_L_bF_buf11), .Y(_416_) );
	AOI21X1 AOI21X1_148 ( .A(_415_), .B(_261__bF_buf4), .C(_416_), .Y(_256__109_) );
	INVX1 INVX1_113 ( .A(bloque_in_110_), .Y(_417_) );
	OAI21X1 OAI21X1_149 ( .A(_261__bF_buf3), .B(RAM_entrada_89_), .C(reset_L_bF_buf10), .Y(_418_) );
	AOI21X1 AOI21X1_149 ( .A(_417_), .B(_261__bF_buf2), .C(_418_), .Y(_256__110_) );
	INVX1 INVX1_114 ( .A(bloque_in_111_), .Y(_419_) );
	OAI21X1 OAI21X1_150 ( .A(_261__bF_buf1), .B(RAM_entrada_88_), .C(reset_L_bF_buf9), .Y(_420_) );
	AOI21X1 AOI21X1_150 ( .A(_419_), .B(_261__bF_buf0), .C(_420_), .Y(_256__111_) );
	INVX1 INVX1_115 ( .A(bloque_in_112_), .Y(_421_) );
	OAI21X1 OAI21X1_151 ( .A(_261__bF_buf15), .B(RAM_entrada_85_), .C(reset_L_bF_buf8), .Y(_422_) );
	AOI21X1 AOI21X1_151 ( .A(_421_), .B(_261__bF_buf14), .C(_422_), .Y(_256__112_) );
	INVX1 INVX1_116 ( .A(bloque_in_113_), .Y(_423_) );
	OAI21X1 OAI21X1_152 ( .A(_261__bF_buf13), .B(RAM_entrada_89_), .C(reset_L_bF_buf7), .Y(_424_) );
	AOI21X1 AOI21X1_152 ( .A(_423_), .B(_261__bF_buf12), .C(_424_), .Y(_256__113_) );
	INVX1 INVX1_117 ( .A(bloque_in_114_), .Y(_425_) );
	OAI21X1 OAI21X1_153 ( .A(_261__bF_buf11), .B(RAM_entrada_82_), .C(reset_L_bF_buf6), .Y(_426_) );
	AOI21X1 AOI21X1_153 ( .A(_425_), .B(_261__bF_buf10), .C(_426_), .Y(_256__114_) );
	INVX1 INVX1_118 ( .A(bloque_in_115_), .Y(_427_) );
	OAI21X1 OAI21X1_154 ( .A(_261__bF_buf9), .B(RAM_entrada_84_), .C(reset_L_bF_buf5), .Y(_428_) );
	AOI21X1 AOI21X1_154 ( .A(_427_), .B(_261__bF_buf8), .C(_428_), .Y(_256__115_) );
	INVX1 INVX1_119 ( .A(bloque_in_116_), .Y(_429_) );
	OAI21X1 OAI21X1_155 ( .A(_261__bF_buf7), .B(RAM_entrada_84_), .C(reset_L_bF_buf4), .Y(_430_) );
	AOI21X1 AOI21X1_155 ( .A(_429_), .B(_261__bF_buf6), .C(_430_), .Y(_256__116_) );
	INVX1 INVX1_120 ( .A(bloque_in_117_), .Y(_431_) );
	OAI21X1 OAI21X1_156 ( .A(_261__bF_buf5), .B(RAM_entrada_85_), .C(reset_L_bF_buf3), .Y(_432_) );
	AOI21X1 AOI21X1_156 ( .A(_431_), .B(_261__bF_buf4), .C(_432_), .Y(_256__117_) );
	INVX1 INVX1_121 ( .A(bloque_in_118_), .Y(_433_) );
	OAI21X1 OAI21X1_157 ( .A(_261__bF_buf3), .B(RAM_entrada_86_), .C(reset_L_bF_buf2), .Y(_434_) );
	AOI21X1 AOI21X1_157 ( .A(_433_), .B(_261__bF_buf2), .C(_434_), .Y(_256__118_) );
	INVX1 INVX1_122 ( .A(bloque_in_119_), .Y(_435_) );
	OAI21X1 OAI21X1_158 ( .A(_261__bF_buf1), .B(gnd), .C(reset_L_bF_buf1), .Y(_436_) );
	AOI21X1 AOI21X1_158 ( .A(_435_), .B(_261__bF_buf0), .C(_436_), .Y(_256__119_) );
	INVX1 INVX1_123 ( .A(bloque_in_120_), .Y(_437_) );
	OAI21X1 OAI21X1_159 ( .A(_261__bF_buf15), .B(RAM_entrada_88_), .C(reset_L_bF_buf0), .Y(_438_) );
	AOI21X1 AOI21X1_159 ( .A(_437_), .B(_261__bF_buf14), .C(_438_), .Y(_256__120_) );
	INVX1 INVX1_124 ( .A(bloque_in_121_), .Y(_439_) );
	OAI21X1 OAI21X1_160 ( .A(_261__bF_buf13), .B(RAM_entrada_89_), .C(reset_L_bF_buf11), .Y(_440_) );
	AOI21X1 AOI21X1_160 ( .A(_439_), .B(_261__bF_buf12), .C(_440_), .Y(_256__121_) );
	INVX1 INVX1_125 ( .A(bloque_in_122_), .Y(_441_) );
	OAI21X1 OAI21X1_161 ( .A(_261__bF_buf11), .B(RAM_entrada_94_), .C(reset_L_bF_buf10), .Y(_442_) );
	AOI21X1 AOI21X1_161 ( .A(_441_), .B(_261__bF_buf10), .C(_442_), .Y(_256__122_) );
	INVX1 INVX1_126 ( .A(bloque_in_123_), .Y(_443_) );
	OAI21X1 OAI21X1_162 ( .A(_261__bF_buf9), .B(vdd), .C(reset_L_bF_buf9), .Y(_444_) );
	AOI21X1 AOI21X1_162 ( .A(_443_), .B(_261__bF_buf8), .C(_444_), .Y(_256__123_) );
	INVX1 INVX1_127 ( .A(bloque_in_124_), .Y(_445_) );
	OAI21X1 OAI21X1_163 ( .A(_261__bF_buf7), .B(RAM_entrada_92_), .C(reset_L_bF_buf8), .Y(_446_) );
	AOI21X1 AOI21X1_163 ( .A(_445_), .B(_261__bF_buf6), .C(_446_), .Y(_256__124_) );
	INVX1 INVX1_128 ( .A(bloque_in_125_), .Y(_447_) );
	OAI21X1 OAI21X1_164 ( .A(_261__bF_buf5), .B(RAM_entrada_93_), .C(reset_L_bF_buf7), .Y(_448_) );
	AOI21X1 AOI21X1_164 ( .A(_447_), .B(_261__bF_buf4), .C(_448_), .Y(_256__125_) );
	INVX1 INVX1_129 ( .A(bloque_in_126_), .Y(_449_) );
	OAI21X1 OAI21X1_165 ( .A(_261__bF_buf3), .B(RAM_entrada_94_), .C(reset_L_bF_buf6), .Y(_450_) );
	AOI21X1 AOI21X1_165 ( .A(_449_), .B(_261__bF_buf2), .C(_450_), .Y(_256__126_) );
	INVX1 INVX1_130 ( .A(bloque_in_127_), .Y(_451_) );
	OAI21X1 OAI21X1_166 ( .A(_261__bF_buf1), .B(RAM_entrada_95_), .C(reset_L_bF_buf5), .Y(_452_) );
	AOI21X1 AOI21X1_166 ( .A(_451_), .B(_261__bF_buf0), .C(_452_), .Y(_256__127_) );
	INVX1 INVX1_131 ( .A(bloque_in_0_), .Y(_453_) );
	OAI21X1 OAI21X1_167 ( .A(_261__bF_buf15), .B(_2__0_), .C(reset_L_bF_buf4), .Y(_454_) );
	AOI21X1 AOI21X1_167 ( .A(_453_), .B(_261__bF_buf14), .C(_454_), .Y(_256__0_) );
	INVX1 INVX1_132 ( .A(bloque_in_1_), .Y(_455_) );
	OAI21X1 OAI21X1_168 ( .A(_261__bF_buf13), .B(_2__1_), .C(reset_L_bF_buf3), .Y(_456_) );
	AOI21X1 AOI21X1_168 ( .A(_455_), .B(_261__bF_buf12), .C(_456_), .Y(_256__1_) );
	INVX1 INVX1_133 ( .A(bloque_in_2_), .Y(_457_) );
	OAI21X1 OAI21X1_169 ( .A(_261__bF_buf11), .B(_2__2_), .C(reset_L_bF_buf2), .Y(_458_) );
	AOI21X1 AOI21X1_169 ( .A(_457_), .B(_261__bF_buf10), .C(_458_), .Y(_256__2_) );
	INVX1 INVX1_134 ( .A(bloque_in_3_), .Y(_459_) );
	OAI21X1 OAI21X1_170 ( .A(_261__bF_buf9), .B(_2__3_), .C(reset_L_bF_buf1), .Y(_460_) );
	AOI21X1 AOI21X1_170 ( .A(_459_), .B(_261__bF_buf8), .C(_460_), .Y(_256__3_) );
	INVX1 INVX1_135 ( .A(bloque_in_4_), .Y(_461_) );
	OAI21X1 OAI21X1_171 ( .A(_261__bF_buf7), .B(_2__4_), .C(reset_L_bF_buf0), .Y(_462_) );
	AOI21X1 AOI21X1_171 ( .A(_461_), .B(_261__bF_buf6), .C(_462_), .Y(_256__4_) );
	INVX1 INVX1_136 ( .A(bloque_in_5_), .Y(_463_) );
	OAI21X1 OAI21X1_172 ( .A(_261__bF_buf5), .B(_2__5_), .C(reset_L_bF_buf11), .Y(_464_) );
	AOI21X1 AOI21X1_172 ( .A(_463_), .B(_261__bF_buf4), .C(_464_), .Y(_256__5_) );
	INVX1 INVX1_137 ( .A(bloque_in_6_), .Y(_465_) );
	OAI21X1 OAI21X1_173 ( .A(_261__bF_buf3), .B(_2__6_), .C(reset_L_bF_buf10), .Y(_466_) );
	AOI21X1 AOI21X1_173 ( .A(_465_), .B(_261__bF_buf2), .C(_466_), .Y(_256__6_) );
	INVX1 INVX1_138 ( .A(bloque_in_7_), .Y(_467_) );
	OAI21X1 OAI21X1_174 ( .A(_261__bF_buf1), .B(_2__7_), .C(reset_L_bF_buf9), .Y(_468_) );
	AOI21X1 AOI21X1_174 ( .A(_467_), .B(_261__bF_buf0), .C(_468_), .Y(_256__7_) );
	INVX1 INVX1_139 ( .A(bloque_in_8_), .Y(_469_) );
	OAI21X1 OAI21X1_175 ( .A(_261__bF_buf15), .B(_2__8_), .C(reset_L_bF_buf8), .Y(_470_) );
	AOI21X1 AOI21X1_175 ( .A(_469_), .B(_261__bF_buf14), .C(_470_), .Y(_256__8_) );
	INVX1 INVX1_140 ( .A(bloque_in_9_), .Y(_471_) );
	OAI21X1 OAI21X1_176 ( .A(_261__bF_buf13), .B(_2__9_), .C(reset_L_bF_buf7), .Y(_472_) );
	AOI21X1 AOI21X1_176 ( .A(_471_), .B(_261__bF_buf12), .C(_472_), .Y(_256__9_) );
	INVX1 INVX1_141 ( .A(bloque_in_10_), .Y(_473_) );
	OAI21X1 OAI21X1_177 ( .A(_261__bF_buf11), .B(_2__10_), .C(reset_L_bF_buf6), .Y(_474_) );
	AOI21X1 AOI21X1_177 ( .A(_473_), .B(_261__bF_buf10), .C(_474_), .Y(_256__10_) );
	INVX1 INVX1_142 ( .A(bloque_in_11_), .Y(_475_) );
	OAI21X1 OAI21X1_178 ( .A(_261__bF_buf9), .B(_2__11_), .C(reset_L_bF_buf5), .Y(_476_) );
	AOI21X1 AOI21X1_178 ( .A(_475_), .B(_261__bF_buf8), .C(_476_), .Y(_256__11_) );
	INVX1 INVX1_143 ( .A(bloque_in_12_), .Y(_477_) );
	OAI21X1 OAI21X1_179 ( .A(_261__bF_buf7), .B(_2__12_), .C(reset_L_bF_buf4), .Y(_478_) );
	AOI21X1 AOI21X1_179 ( .A(_477_), .B(_261__bF_buf6), .C(_478_), .Y(_256__12_) );
	INVX1 INVX1_144 ( .A(bloque_in_13_), .Y(_479_) );
	OAI21X1 OAI21X1_180 ( .A(_261__bF_buf5), .B(_2__13_), .C(reset_L_bF_buf3), .Y(_480_) );
	AOI21X1 AOI21X1_180 ( .A(_479_), .B(_261__bF_buf4), .C(_480_), .Y(_256__13_) );
	INVX1 INVX1_145 ( .A(bloque_in_14_), .Y(_481_) );
	OAI21X1 OAI21X1_181 ( .A(_261__bF_buf3), .B(_2__14_), .C(reset_L_bF_buf2), .Y(_482_) );
	AOI21X1 AOI21X1_181 ( .A(_481_), .B(_261__bF_buf2), .C(_482_), .Y(_256__14_) );
	INVX1 INVX1_146 ( .A(bloque_in_15_), .Y(_483_) );
	OAI21X1 OAI21X1_182 ( .A(_261__bF_buf1), .B(_2__15_), .C(reset_L_bF_buf1), .Y(_484_) );
	AOI21X1 AOI21X1_182 ( .A(_483_), .B(_261__bF_buf0), .C(_484_), .Y(_256__15_) );
	INVX1 INVX1_147 ( .A(bloque_in_16_), .Y(_485_) );
	OAI21X1 OAI21X1_183 ( .A(_261__bF_buf15), .B(_2__16_), .C(reset_L_bF_buf0), .Y(_486_) );
	AOI21X1 AOI21X1_183 ( .A(_485_), .B(_261__bF_buf14), .C(_486_), .Y(_256__16_) );
	INVX1 INVX1_148 ( .A(bloque_in_17_), .Y(_487_) );
	OAI21X1 OAI21X1_184 ( .A(_261__bF_buf13), .B(_2__17_), .C(reset_L_bF_buf11), .Y(_488_) );
	AOI21X1 AOI21X1_184 ( .A(_487_), .B(_261__bF_buf12), .C(_488_), .Y(_256__17_) );
	INVX1 INVX1_149 ( .A(bloque_in_18_), .Y(_489_) );
	OAI21X1 OAI21X1_185 ( .A(_261__bF_buf11), .B(_2__18_), .C(reset_L_bF_buf10), .Y(_490_) );
	AOI21X1 AOI21X1_185 ( .A(_489_), .B(_261__bF_buf10), .C(_490_), .Y(_256__18_) );
	INVX1 INVX1_150 ( .A(bloque_in_19_), .Y(_491_) );
	OAI21X1 OAI21X1_186 ( .A(_261__bF_buf9), .B(_2__19_), .C(reset_L_bF_buf9), .Y(_492_) );
	AOI21X1 AOI21X1_186 ( .A(_491_), .B(_261__bF_buf8), .C(_492_), .Y(_256__19_) );
	INVX1 INVX1_151 ( .A(bloque_in_20_), .Y(_493_) );
	OAI21X1 OAI21X1_187 ( .A(_261__bF_buf7), .B(_2__20_), .C(reset_L_bF_buf8), .Y(_494_) );
	AOI21X1 AOI21X1_187 ( .A(_493_), .B(_261__bF_buf6), .C(_494_), .Y(_256__20_) );
	INVX1 INVX1_152 ( .A(bloque_in_21_), .Y(_495_) );
	OAI21X1 OAI21X1_188 ( .A(_261__bF_buf5), .B(_2__21_), .C(reset_L_bF_buf7), .Y(_496_) );
	AOI21X1 AOI21X1_188 ( .A(_495_), .B(_261__bF_buf4), .C(_496_), .Y(_256__21_) );
	INVX1 INVX1_153 ( .A(bloque_in_22_), .Y(_497_) );
	OAI21X1 OAI21X1_189 ( .A(_261__bF_buf3), .B(_2__22_), .C(reset_L_bF_buf6), .Y(_498_) );
	AOI21X1 AOI21X1_189 ( .A(_497_), .B(_261__bF_buf2), .C(_498_), .Y(_256__22_) );
	INVX1 INVX1_154 ( .A(bloque_in_23_), .Y(_499_) );
	OAI21X1 OAI21X1_190 ( .A(_261__bF_buf1), .B(_2__23_), .C(reset_L_bF_buf5), .Y(_500_) );
	AOI21X1 AOI21X1_190 ( .A(_499_), .B(_261__bF_buf0), .C(_500_), .Y(_256__23_) );
	INVX1 INVX1_155 ( .A(bloque_in_24_), .Y(_501_) );
	OAI21X1 OAI21X1_191 ( .A(_261__bF_buf15), .B(_2__24_), .C(reset_L_bF_buf4), .Y(_502_) );
	AOI21X1 AOI21X1_191 ( .A(_501_), .B(_261__bF_buf14), .C(_502_), .Y(_256__24_) );
	INVX1 INVX1_156 ( .A(bloque_in_25_), .Y(_503_) );
	OAI21X1 OAI21X1_192 ( .A(_261__bF_buf13), .B(_2__25_), .C(reset_L_bF_buf3), .Y(_504_) );
	AOI21X1 AOI21X1_192 ( .A(_503_), .B(_261__bF_buf12), .C(_504_), .Y(_256__25_) );
	INVX1 INVX1_157 ( .A(bloque_in_26_), .Y(_505_) );
	OAI21X1 OAI21X1_193 ( .A(_261__bF_buf11), .B(_2__26_), .C(reset_L_bF_buf2), .Y(_506_) );
	AOI21X1 AOI21X1_193 ( .A(_505_), .B(_261__bF_buf10), .C(_506_), .Y(_256__26_) );
	INVX1 INVX1_158 ( .A(bloque_in_27_), .Y(_507_) );
	OAI21X1 OAI21X1_194 ( .A(_261__bF_buf9), .B(_2__27_), .C(reset_L_bF_buf1), .Y(_508_) );
	AOI21X1 AOI21X1_194 ( .A(_507_), .B(_261__bF_buf8), .C(_508_), .Y(_256__27_) );
	INVX1 INVX1_159 ( .A(bloque_in_28_), .Y(_509_) );
	OAI21X1 OAI21X1_195 ( .A(_261__bF_buf7), .B(_2__28_), .C(reset_L_bF_buf0), .Y(_510_) );
	AOI21X1 AOI21X1_195 ( .A(_509_), .B(_261__bF_buf6), .C(_510_), .Y(_256__28_) );
	INVX1 INVX1_160 ( .A(bloque_in_29_), .Y(_511_) );
	OAI21X1 OAI21X1_196 ( .A(_261__bF_buf5), .B(_2__29_), .C(reset_L_bF_buf11), .Y(_512_) );
	AOI21X1 AOI21X1_196 ( .A(_511_), .B(_261__bF_buf4), .C(_512_), .Y(_256__29_) );
	INVX1 INVX1_161 ( .A(bloque_in_30_), .Y(_513_) );
	OAI21X1 OAI21X1_197 ( .A(_261__bF_buf3), .B(_2__30_), .C(reset_L_bF_buf10), .Y(_514_) );
	AOI21X1 AOI21X1_197 ( .A(_513_), .B(_261__bF_buf2), .C(_514_), .Y(_256__30_) );
	INVX1 INVX1_162 ( .A(bloque_in_31_), .Y(_515_) );
	OAI21X1 OAI21X1_198 ( .A(_261__bF_buf1), .B(_2__31_), .C(reset_L_bF_buf9), .Y(_516_) );
	AOI21X1 AOI21X1_198 ( .A(_515_), .B(_261__bF_buf0), .C(_516_), .Y(_256__31_) );
	DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf5), .D(_256__0_), .Q(bloque_in_0_) );
	DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf4), .D(_256__1_), .Q(bloque_in_1_) );
	DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf3), .D(_256__2_), .Q(bloque_in_2_) );
	DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf2), .D(_256__3_), .Q(bloque_in_3_) );
	DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf1), .D(_256__4_), .Q(bloque_in_4_) );
	DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf0), .D(_256__5_), .Q(bloque_in_5_) );
	DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf76), .D(_256__6_), .Q(bloque_in_6_) );
	DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf75), .D(_256__7_), .Q(bloque_in_7_) );
	DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf74), .D(_256__8_), .Q(bloque_in_8_) );
	DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf73), .D(_256__9_), .Q(bloque_in_9_) );
	DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf72), .D(_256__10_), .Q(bloque_in_10_) );
	DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf71), .D(_256__11_), .Q(bloque_in_11_) );
	DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf70), .D(_256__12_), .Q(bloque_in_12_) );
	DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf69), .D(_256__13_), .Q(bloque_in_13_) );
	DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf68), .D(_256__14_), .Q(bloque_in_14_) );
	DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf67), .D(_256__15_), .Q(bloque_in_15_) );
	DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf66), .D(_256__16_), .Q(bloque_in_16_) );
	DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf65), .D(_256__17_), .Q(bloque_in_17_) );
	DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf64), .D(_256__18_), .Q(bloque_in_18_) );
	DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf63), .D(_256__19_), .Q(bloque_in_19_) );
	DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf62), .D(_256__20_), .Q(bloque_in_20_) );
	DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf61), .D(_256__21_), .Q(bloque_in_21_) );
	DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf60), .D(_256__22_), .Q(bloque_in_22_) );
	DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf59), .D(_256__23_), .Q(bloque_in_23_) );
	DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf58), .D(_256__24_), .Q(bloque_in_24_) );
	DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf57), .D(_256__25_), .Q(bloque_in_25_) );
	DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf56), .D(_256__26_), .Q(bloque_in_26_) );
	DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf55), .D(_256__27_), .Q(bloque_in_27_) );
	DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf54), .D(_256__28_), .Q(bloque_in_28_) );
	DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf53), .D(_256__29_), .Q(bloque_in_29_) );
	DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf52), .D(_256__30_), .Q(bloque_in_30_) );
	DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf51), .D(_256__31_), .Q(bloque_in_31_) );
	DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf50), .D(_256__32_), .Q(bloque_in_32_) );
	DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf49), .D(_256__33_), .Q(bloque_in_33_) );
	DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf48), .D(_256__34_), .Q(bloque_in_34_) );
	DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf47), .D(_256__35_), .Q(bloque_in_35_) );
	DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf46), .D(_256__36_), .Q(bloque_in_36_) );
	DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf45), .D(_256__37_), .Q(bloque_in_37_) );
	DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf44), .D(_256__38_), .Q(bloque_in_38_) );
	DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf43), .D(_256__39_), .Q(bloque_in_39_) );
	DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf42), .D(_256__40_), .Q(bloque_in_40_) );
	DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf41), .D(_256__41_), .Q(bloque_in_41_) );
	DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf40), .D(_256__42_), .Q(bloque_in_42_) );
	DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf39), .D(_256__43_), .Q(bloque_in_43_) );
	DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf38), .D(_256__44_), .Q(bloque_in_44_) );
	DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf37), .D(_256__45_), .Q(bloque_in_45_) );
	DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf36), .D(_256__46_), .Q(bloque_in_46_) );
	DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf35), .D(_256__47_), .Q(bloque_in_47_) );
	DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf34), .D(_256__48_), .Q(bloque_in_48_) );
	DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf33), .D(_256__49_), .Q(bloque_in_49_) );
	DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf32), .D(_256__50_), .Q(bloque_in_50_) );
	DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf31), .D(_256__51_), .Q(bloque_in_51_) );
	DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf30), .D(_256__52_), .Q(bloque_in_52_) );
	DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf29), .D(_256__53_), .Q(bloque_in_53_) );
	DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf28), .D(_256__54_), .Q(bloque_in_54_) );
	DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf27), .D(_256__55_), .Q(bloque_in_55_) );
	DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf26), .D(_256__56_), .Q(bloque_in_56_) );
	DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf25), .D(_256__57_), .Q(bloque_in_57_) );
	DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf24), .D(_256__58_), .Q(bloque_in_58_) );
	DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf23), .D(_256__59_), .Q(bloque_in_59_) );
	DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf22), .D(_256__60_), .Q(bloque_in_60_) );
	DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf21), .D(_256__61_), .Q(bloque_in_61_) );
	DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf20), .D(_256__62_), .Q(bloque_in_62_) );
	DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf19), .D(_256__63_), .Q(bloque_in_63_) );
	DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf18), .D(_256__64_), .Q(bloque_in_64_) );
	DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf17), .D(_256__65_), .Q(bloque_in_65_) );
	DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf16), .D(_256__66_), .Q(bloque_in_66_) );
	DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf15), .D(_256__67_), .Q(bloque_in_67_) );
	DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf14), .D(_256__68_), .Q(bloque_in_68_) );
	DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf13), .D(_256__69_), .Q(bloque_in_69_) );
	DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf12), .D(_256__70_), .Q(bloque_in_70_) );
	DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf11), .D(_256__71_), .Q(bloque_in_71_) );
	DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf10), .D(_256__72_), .Q(bloque_in_72_) );
	DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf9), .D(_256__73_), .Q(bloque_in_73_) );
	DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf8), .D(_256__74_), .Q(bloque_in_74_) );
	DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf7), .D(_256__75_), .Q(bloque_in_75_) );
	DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf6), .D(_256__76_), .Q(bloque_in_76_) );
	DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf5), .D(_256__77_), .Q(bloque_in_77_) );
	DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf4), .D(_256__78_), .Q(bloque_in_78_) );
	DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf3), .D(_256__79_), .Q(bloque_in_79_) );
	DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf2), .D(_256__80_), .Q(bloque_in_80_) );
	DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf1), .D(_256__81_), .Q(bloque_in_81_) );
	DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf0), .D(_256__82_), .Q(bloque_in_82_) );
	DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf76), .D(_256__83_), .Q(bloque_in_83_) );
	DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf75), .D(_256__84_), .Q(bloque_in_84_) );
	DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf74), .D(_256__85_), .Q(bloque_in_85_) );
	DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf73), .D(_256__86_), .Q(bloque_in_86_) );
	DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf72), .D(_256__87_), .Q(bloque_in_87_) );
	DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf71), .D(_256__88_), .Q(bloque_in_88_) );
	DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf70), .D(_256__89_), .Q(bloque_in_89_) );
	DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf69), .D(_256__90_), .Q(bloque_in_90_) );
	DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf68), .D(_256__91_), .Q(bloque_in_91_) );
	DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf67), .D(_256__92_), .Q(bloque_in_92_) );
	DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf66), .D(_256__93_), .Q(bloque_in_93_) );
	DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf65), .D(_256__94_), .Q(bloque_in_94_) );
	DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf64), .D(_256__95_), .Q(bloque_in_95_) );
	DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf63), .D(_256__96_), .Q(bloque_in_96_) );
	DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf62), .D(_256__97_), .Q(bloque_in_97_) );
	DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf61), .D(_256__98_), .Q(bloque_in_98_) );
	DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf60), .D(_256__99_), .Q(bloque_in_99_) );
	DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf59), .D(_256__100_), .Q(bloque_in_100_) );
	DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf58), .D(_256__101_), .Q(bloque_in_101_) );
	DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf57), .D(_256__102_), .Q(bloque_in_102_) );
	DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf56), .D(_256__103_), .Q(bloque_in_103_) );
	DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf55), .D(_256__104_), .Q(bloque_in_104_) );
	DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf54), .D(_256__105_), .Q(bloque_in_105_) );
	DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf53), .D(_256__106_), .Q(bloque_in_106_) );
	DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf52), .D(_256__107_), .Q(bloque_in_107_) );
	DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf51), .D(_256__108_), .Q(bloque_in_108_) );
	DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf50), .D(_256__109_), .Q(bloque_in_109_) );
	DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf49), .D(_256__110_), .Q(bloque_in_110_) );
	DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf48), .D(_256__111_), .Q(bloque_in_111_) );
	DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf47), .D(_256__112_), .Q(bloque_in_112_) );
	DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf46), .D(_256__113_), .Q(bloque_in_113_) );
	DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf45), .D(_256__114_), .Q(bloque_in_114_) );
	DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf44), .D(_256__115_), .Q(bloque_in_115_) );
	DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf43), .D(_256__116_), .Q(bloque_in_116_) );
	DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf42), .D(_256__117_), .Q(bloque_in_117_) );
	DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf41), .D(_256__118_), .Q(bloque_in_118_) );
	DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf40), .D(_256__119_), .Q(bloque_in_119_) );
	DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf39), .D(_256__120_), .Q(bloque_in_120_) );
	DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf38), .D(_256__121_), .Q(bloque_in_121_) );
	DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf37), .D(_256__122_), .Q(bloque_in_122_) );
	DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf36), .D(_256__123_), .Q(bloque_in_123_) );
	DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf35), .D(_256__124_), .Q(bloque_in_124_) );
	DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf34), .D(_256__125_), .Q(bloque_in_125_) );
	DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf33), .D(_256__126_), .Q(bloque_in_126_) );
	DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf32), .D(_256__127_), .Q(bloque_in_127_) );
	NOR2X1 NOR2X1_25 ( .A(reset_L_bF_buf8), .B(_1__bF_buf1), .Y(_519_) );
	INVX2 INVX2_1 ( .A(_519_), .Y(_520_) );
	AND2X2 AND2X2_2 ( .A(_520_), .B(gen_nonce_synth_rand_0_), .Y(_518__0_) );
	OR2X2 OR2X2_6 ( .A(_519_), .B(gen_nonce_synth_rand_1_), .Y(_518__1_) );
	INVX1 INVX1_163 ( .A(gen_nonce_synth_rand_2_), .Y(_521_) );
	NOR2X1 NOR2X1_26 ( .A(_521_), .B(_519_), .Y(_518__2_) );
	INVX1 INVX1_164 ( .A(gen_nonce_synth_rand_3_), .Y(_522_) );
	OAI21X1 OAI21X1_199 ( .A(reset_L_bF_buf7), .B(_1__bF_buf0), .C(_522_), .Y(_518__3_) );
	AND2X2 AND2X2_3 ( .A(_520_), .B(gen_nonce_synth_rand_4_), .Y(_518__4_) );
	AND2X2 AND2X2_4 ( .A(_520_), .B(gen_nonce_synth_rand_5_), .Y(_518__5_) );
	INVX1 INVX1_165 ( .A(gen_nonce_synth_rand_6_), .Y(_523_) );
	OAI21X1 OAI21X1_200 ( .A(reset_L_bF_buf6), .B(_1__bF_buf5), .C(_523_), .Y(_518__6_) );
	AND2X2 AND2X2_5 ( .A(_520_), .B(gen_nonce_synth_rand_7_), .Y(_518__7_) );
	INVX1 INVX1_166 ( .A(gen_nonce_synth_rand_8_), .Y(_524_) );
	NOR2X1 NOR2X1_27 ( .A(_524_), .B(_519_), .Y(_518__8_) );
	INVX1 INVX1_167 ( .A(gen_nonce_synth_rand_9_), .Y(_525_) );
	OAI21X1 OAI21X1_201 ( .A(reset_L_bF_buf5), .B(_1__bF_buf4), .C(_525_), .Y(_518__9_) );
	INVX1 INVX1_168 ( .A(gen_nonce_synth_rand_10_), .Y(_526_) );
	NOR2X1 NOR2X1_28 ( .A(_526_), .B(_519_), .Y(_518__10_) );
	INVX1 INVX1_169 ( .A(gen_nonce_synth_rand_11_), .Y(_527_) );
	NOR2X1 NOR2X1_29 ( .A(_527_), .B(_519_), .Y(_518__11_) );
	INVX1 INVX1_170 ( .A(gen_nonce_synth_rand_12_), .Y(_528_) );
	OAI21X1 OAI21X1_202 ( .A(reset_L_bF_buf4), .B(_1__bF_buf3), .C(_528_), .Y(_518__12_) );
	INVX1 INVX1_171 ( .A(gen_nonce_synth_rand_13_), .Y(_529_) );
	OAI21X1 OAI21X1_203 ( .A(reset_L_bF_buf3), .B(_1__bF_buf2), .C(_529_), .Y(_518__13_) );
	INVX1 INVX1_172 ( .A(gen_nonce_synth_rand_14_), .Y(_530_) );
	OAI21X1 OAI21X1_204 ( .A(reset_L_bF_buf2), .B(_1__bF_buf1), .C(_530_), .Y(_518__14_) );
	INVX1 INVX1_173 ( .A(gen_nonce_synth_rand_15_), .Y(_531_) );
	NOR2X1 NOR2X1_30 ( .A(_531_), .B(_519_), .Y(_518__15_) );
	INVX1 INVX1_174 ( .A(gen_nonce_synth_rand_16_), .Y(_532_) );
	OAI21X1 OAI21X1_205 ( .A(reset_L_bF_buf1), .B(_1__bF_buf0), .C(_532_), .Y(_518__16_) );
	INVX1 INVX1_175 ( .A(gen_nonce_synth_rand_17_), .Y(_533_) );
	OAI21X1 OAI21X1_206 ( .A(reset_L_bF_buf0), .B(_1__bF_buf5), .C(_533_), .Y(_518__17_) );
	INVX1 INVX1_176 ( .A(gen_nonce_synth_rand_18_), .Y(_534_) );
	NOR2X1 NOR2X1_31 ( .A(_534_), .B(_519_), .Y(_518__18_) );
	INVX1 INVX1_177 ( .A(gen_nonce_synth_rand_19_), .Y(_535_) );
	OAI21X1 OAI21X1_207 ( .A(reset_L_bF_buf11), .B(_1__bF_buf4), .C(_535_), .Y(_518__19_) );
	INVX1 INVX1_178 ( .A(gen_nonce_synth_rand_20_), .Y(_536_) );
	NOR2X1 NOR2X1_32 ( .A(_536_), .B(_519_), .Y(_518__20_) );
	INVX1 INVX1_179 ( .A(gen_nonce_synth_rand_21_), .Y(_537_) );
	NOR2X1 NOR2X1_33 ( .A(_537_), .B(_519_), .Y(_518__21_) );
	INVX1 INVX1_180 ( .A(gen_nonce_synth_rand_22_), .Y(_538_) );
	OAI21X1 OAI21X1_208 ( .A(reset_L_bF_buf10), .B(_1__bF_buf3), .C(_538_), .Y(_518__22_) );
	INVX1 INVX1_181 ( .A(gen_nonce_synth_rand_23_), .Y(_539_) );
	NOR2X1 NOR2X1_34 ( .A(_539_), .B(_519_), .Y(_518__23_) );
	INVX1 INVX1_182 ( .A(gen_nonce_synth_rand_24_), .Y(_540_) );
	OAI21X1 OAI21X1_209 ( .A(reset_L_bF_buf9), .B(_1__bF_buf2), .C(_540_), .Y(_518__24_) );
	INVX1 INVX1_183 ( .A(gen_nonce_synth_rand_25_), .Y(_541_) );
	OAI21X1 OAI21X1_210 ( .A(reset_L_bF_buf8), .B(_1__bF_buf1), .C(_541_), .Y(_518__25_) );
	AND2X2 AND2X2_6 ( .A(_520_), .B(gen_nonce_synth_rand_26_), .Y(_518__26_) );
	AND2X2 AND2X2_7 ( .A(_520_), .B(gen_nonce_synth_rand_27_), .Y(_518__27_) );
	INVX1 INVX1_184 ( .A(gen_nonce_synth_rand_28_), .Y(_542_) );
	NOR2X1 NOR2X1_35 ( .A(_542_), .B(_519_), .Y(_518__28_) );
	INVX1 INVX1_185 ( .A(gen_nonce_synth_rand_29_), .Y(_543_) );
	OAI21X1 OAI21X1_211 ( .A(reset_L_bF_buf7), .B(_1__bF_buf0), .C(_543_), .Y(_518__29_) );
	AND2X2 AND2X2_8 ( .A(_520_), .B(gen_nonce_synth_rand_30_), .Y(_518__30_) );
	AND2X2 AND2X2_9 ( .A(_520_), .B(gen_nonce_synth_rand_31_), .Y(_518__31_) );
	INVX4 INVX4_1 ( .A(_1__bF_buf5), .Y(_544_) );
	INVX8 INVX8_2 ( .A(comparador_valid_bF_buf4), .Y(_545_) );
	NAND3X1 NAND3X1_62 ( .A(gen_nonce_synth_rand_0_), .B(_544_), .C(_545__bF_buf4), .Y(_546_) );
	AND2X2 AND2X2_10 ( .A(_546_), .B(_2__0_), .Y(_547_) );
	OAI21X1 OAI21X1_212 ( .A(_546_), .B(_2__0_), .C(_520_), .Y(_548_) );
	OR2X2 OR2X2_7 ( .A(_547_), .B(_548_), .Y(_517__0_) );
	INVX1 INVX1_186 ( .A(_2__1_), .Y(_549_) );
	NAND2X1 NAND2X1_38 ( .A(gen_nonce_synth_rand_0_), .B(_2__0_), .Y(_550_) );
	AND2X2 AND2X2_11 ( .A(gen_nonce_synth_rand_1_), .B(_2__1_), .Y(_551_) );
	NOR2X1 NOR2X1_36 ( .A(gen_nonce_synth_rand_1_), .B(_2__1_), .Y(_552_) );
	NOR2X1 NOR2X1_37 ( .A(_552_), .B(_551_), .Y(_553_) );
	XNOR2X1 XNOR2X1_1 ( .A(_553_), .B(_550_), .Y(_554_) );
	NAND2X1 NAND2X1_39 ( .A(comparador_valid_bF_buf3), .B(_549_), .Y(_555_) );
	OAI21X1 OAI21X1_213 ( .A(_554_), .B(comparador_valid_bF_buf2), .C(_555_), .Y(_556_) );
	NAND2X1 NAND2X1_40 ( .A(reset_L_bF_buf6), .B(_544_), .Y(_557_) );
	INVX4 INVX4_2 ( .A(_557_), .Y(_558_) );
	AOI22X1 AOI22X1_11 ( .A(_1__bF_buf4), .B(_549_), .C(_556_), .D(_558__bF_buf3), .Y(_517__1_) );
	INVX1 INVX1_187 ( .A(_2__2_), .Y(_559_) );
	AND2X2 AND2X2_12 ( .A(gen_nonce_synth_rand_0_), .B(_2__0_), .Y(_560_) );
	OR2X2 OR2X2_8 ( .A(gen_nonce_synth_rand_1_), .B(_2__1_), .Y(_561_) );
	AOI21X1 AOI21X1_199 ( .A(_560_), .B(_561_), .C(_551_), .Y(_562_) );
	XNOR2X1 XNOR2X1_2 ( .A(gen_nonce_synth_rand_2_), .B(_2__2_), .Y(_563_) );
	NOR2X1 NOR2X1_38 ( .A(_563_), .B(_562_), .Y(_564_) );
	AND2X2 AND2X2_13 ( .A(_562_), .B(_563_), .Y(_565_) );
	OAI21X1 OAI21X1_214 ( .A(_565_), .B(_564_), .C(_545__bF_buf3), .Y(_566_) );
	OAI21X1 OAI21X1_215 ( .A(_545__bF_buf2), .B(_2__2_), .C(_566_), .Y(_567_) );
	AOI22X1 AOI22X1_12 ( .A(_1__bF_buf3), .B(_559_), .C(_567_), .D(_558__bF_buf2), .Y(_517__2_) );
	INVX1 INVX1_188 ( .A(_2__3_), .Y(_568_) );
	XNOR2X1 XNOR2X1_3 ( .A(gen_nonce_synth_rand_3_), .B(_2__3_), .Y(_569_) );
	NAND2X1 NAND2X1_41 ( .A(gen_nonce_synth_rand_2_), .B(_2__2_), .Y(_570_) );
	OAI21X1 OAI21X1_216 ( .A(_562_), .B(_563_), .C(_570_), .Y(_571_) );
	OAI21X1 OAI21X1_217 ( .A(_571_), .B(_569_), .C(_545__bF_buf1), .Y(_572_) );
	AOI21X1 AOI21X1_200 ( .A(_569_), .B(_571_), .C(_572_), .Y(_573_) );
	OAI21X1 OAI21X1_218 ( .A(_545__bF_buf0), .B(_2__3_), .C(_558__bF_buf1), .Y(_574_) );
	OAI22X1 OAI22X1_11 ( .A(_544_), .B(_568_), .C(_573_), .D(_574_), .Y(_517__3_) );
	NAND2X1 NAND2X1_42 ( .A(_1__bF_buf2), .B(_2__4_), .Y(_575_) );
	INVX1 INVX1_189 ( .A(_551_), .Y(_576_) );
	OAI21X1 OAI21X1_219 ( .A(_552_), .B(_550_), .C(_576_), .Y(_577_) );
	NAND2X1 NAND2X1_43 ( .A(gen_nonce_synth_rand_2_), .B(_559_), .Y(_578_) );
	NAND2X1 NAND2X1_44 ( .A(_2__2_), .B(_521_), .Y(_579_) );
	NAND2X1 NAND2X1_45 ( .A(gen_nonce_synth_rand_3_), .B(_568_), .Y(_580_) );
	NAND2X1 NAND2X1_46 ( .A(_2__3_), .B(_522_), .Y(_581_) );
	AOI22X1 AOI22X1_13 ( .A(_578_), .B(_579_), .C(_580_), .D(_581_), .Y(_582_) );
	NAND2X1 NAND2X1_47 ( .A(gen_nonce_synth_rand_3_), .B(_2__3_), .Y(_583_) );
	NOR2X1 NOR2X1_39 ( .A(gen_nonce_synth_rand_3_), .B(_2__3_), .Y(_584_) );
	OAI21X1 OAI21X1_220 ( .A(_584_), .B(_570_), .C(_583_), .Y(_585_) );
	AOI21X1 AOI21X1_201 ( .A(_577_), .B(_582_), .C(_585_), .Y(_586_) );
	XNOR2X1 XNOR2X1_4 ( .A(gen_nonce_synth_rand_4_), .B(_2__4_), .Y(_587_) );
	NAND2X1 NAND2X1_48 ( .A(_587_), .B(_586_), .Y(_588_) );
	NOR3X1 NOR3X1_1 ( .A(_563_), .B(_569_), .C(_562_), .Y(_589_) );
	XOR2X1 XOR2X1_1 ( .A(gen_nonce_synth_rand_4_), .B(_2__4_), .Y(_590_) );
	OAI21X1 OAI21X1_221 ( .A(_589_), .B(_585_), .C(_590_), .Y(_591_) );
	AOI21X1 AOI21X1_202 ( .A(_588_), .B(_591_), .C(comparador_valid_bF_buf1), .Y(_592_) );
	OAI21X1 OAI21X1_222 ( .A(_545__bF_buf4), .B(_2__4_), .C(_558__bF_buf0), .Y(_593_) );
	OAI21X1 OAI21X1_223 ( .A(_592_), .B(_593_), .C(_575_), .Y(_517__4_) );
	NAND2X1 NAND2X1_49 ( .A(gen_nonce_synth_rand_4_), .B(_2__4_), .Y(_594_) );
	OAI21X1 OAI21X1_224 ( .A(_586_), .B(_587_), .C(_594_), .Y(_595_) );
	INVX1 INVX1_190 ( .A(_595_), .Y(_596_) );
	XNOR2X1 XNOR2X1_5 ( .A(gen_nonce_synth_rand_5_), .B(_2__5_), .Y(_597_) );
	AOI21X1 AOI21X1_203 ( .A(_597_), .B(_596_), .C(comparador_valid_bF_buf0), .Y(_598_) );
	OAI21X1 OAI21X1_225 ( .A(_596_), .B(_597_), .C(_598_), .Y(_599_) );
	AOI21X1 AOI21X1_204 ( .A(comparador_valid_bF_buf5), .B(_2__5_), .C(_557_), .Y(_600_) );
	NOR2X1 NOR2X1_40 ( .A(_2__5_), .B(_544_), .Y(_601_) );
	AOI21X1 AOI21X1_205 ( .A(_600_), .B(_599_), .C(_601_), .Y(_517__5_) );
	INVX1 INVX1_191 ( .A(_2__6_), .Y(_602_) );
	NAND2X1 NAND2X1_50 ( .A(gen_nonce_synth_rand_5_), .B(_2__5_), .Y(_603_) );
	NOR2X1 NOR2X1_41 ( .A(gen_nonce_synth_rand_5_), .B(_2__5_), .Y(_604_) );
	OAI21X1 OAI21X1_226 ( .A(_604_), .B(_594_), .C(_603_), .Y(_605_) );
	INVX1 INVX1_192 ( .A(_605_), .Y(_606_) );
	XOR2X1 XOR2X1_2 ( .A(gen_nonce_synth_rand_5_), .B(_2__5_), .Y(_607_) );
	NAND2X1 NAND2X1_51 ( .A(_590_), .B(_607_), .Y(_608_) );
	OAI21X1 OAI21X1_227 ( .A(_586_), .B(_608_), .C(_606_), .Y(_609_) );
	INVX1 INVX1_193 ( .A(_609_), .Y(_610_) );
	XNOR2X1 XNOR2X1_6 ( .A(gen_nonce_synth_rand_6_), .B(_2__6_), .Y(_611_) );
	AOI21X1 AOI21X1_206 ( .A(_611_), .B(_610_), .C(comparador_valid_bF_buf4), .Y(_612_) );
	OAI21X1 OAI21X1_228 ( .A(_610_), .B(_611_), .C(_612_), .Y(_613_) );
	AOI21X1 AOI21X1_207 ( .A(comparador_valid_bF_buf3), .B(_2__6_), .C(_557_), .Y(_614_) );
	AOI22X1 AOI22X1_14 ( .A(_1__bF_buf1), .B(_602_), .C(_613_), .D(_614_), .Y(_517__6_) );
	NAND2X1 NAND2X1_52 ( .A(gen_nonce_synth_rand_6_), .B(_2__6_), .Y(_615_) );
	OAI21X1 OAI21X1_229 ( .A(_610_), .B(_611_), .C(_615_), .Y(_616_) );
	XOR2X1 XOR2X1_3 ( .A(gen_nonce_synth_rand_7_), .B(_2__7_), .Y(_617_) );
	AND2X2 AND2X2_14 ( .A(_616_), .B(_617_), .Y(_618_) );
	OAI21X1 OAI21X1_230 ( .A(_616_), .B(_617_), .C(_545__bF_buf3), .Y(_619_) );
	AOI21X1 AOI21X1_208 ( .A(comparador_valid_bF_buf2), .B(_2__7_), .C(_557_), .Y(_620_) );
	OAI21X1 OAI21X1_231 ( .A(_618_), .B(_619_), .C(_620_), .Y(_621_) );
	OR2X2 OR2X2_9 ( .A(_544_), .B(_2__7_), .Y(_622_) );
	AND2X2 AND2X2_15 ( .A(_621_), .B(_622_), .Y(_517__7_) );
	INVX1 INVX1_194 ( .A(_2__8_), .Y(_623_) );
	NOR2X1 NOR2X1_42 ( .A(_587_), .B(_597_), .Y(_624_) );
	XNOR2X1 XNOR2X1_7 ( .A(gen_nonce_synth_rand_7_), .B(_2__7_), .Y(_625_) );
	NOR2X1 NOR2X1_43 ( .A(_611_), .B(_625_), .Y(_626_) );
	NAND2X1 NAND2X1_53 ( .A(_624_), .B(_626_), .Y(_627_) );
	NAND2X1 NAND2X1_54 ( .A(gen_nonce_synth_rand_7_), .B(_2__7_), .Y(_628_) );
	OAI21X1 OAI21X1_232 ( .A(_625_), .B(_615_), .C(_628_), .Y(_629_) );
	AOI21X1 AOI21X1_209 ( .A(_605_), .B(_626_), .C(_629_), .Y(_630_) );
	OAI21X1 OAI21X1_233 ( .A(_627_), .B(_586_), .C(_630_), .Y(_631_) );
	XOR2X1 XOR2X1_4 ( .A(gen_nonce_synth_rand_8_), .B(_2__8_), .Y(_632_) );
	NAND2X1 NAND2X1_55 ( .A(_632_), .B(_631_), .Y(_633_) );
	OR2X2 OR2X2_10 ( .A(_631_), .B(_632_), .Y(_634_) );
	NAND3X1 NAND3X1_63 ( .A(_545__bF_buf2), .B(_633_), .C(_634_), .Y(_635_) );
	AOI21X1 AOI21X1_210 ( .A(comparador_valid_bF_buf1), .B(_2__8_), .C(_557_), .Y(_636_) );
	AOI22X1 AOI22X1_15 ( .A(_1__bF_buf0), .B(_623_), .C(_635_), .D(_636_), .Y(_517__8_) );
	INVX1 INVX1_195 ( .A(_2__9_), .Y(_637_) );
	XOR2X1 XOR2X1_5 ( .A(gen_nonce_synth_rand_9_), .B(_2__9_), .Y(_638_) );
	INVX1 INVX1_196 ( .A(_638_), .Y(_639_) );
	OAI21X1 OAI21X1_234 ( .A(_524_), .B(_623_), .C(_633_), .Y(_640_) );
	OAI21X1 OAI21X1_235 ( .A(_640_), .B(_639_), .C(_545__bF_buf1), .Y(_641_) );
	AOI21X1 AOI21X1_211 ( .A(_639_), .B(_640_), .C(_641_), .Y(_642_) );
	OAI21X1 OAI21X1_236 ( .A(_545__bF_buf0), .B(_2__9_), .C(_558__bF_buf3), .Y(_643_) );
	OAI22X1 OAI22X1_12 ( .A(_544_), .B(_637_), .C(_642_), .D(_643_), .Y(_517__9_) );
	INVX1 INVX1_197 ( .A(_2__10_), .Y(_644_) );
	NOR2X1 NOR2X1_44 ( .A(_524_), .B(_623_), .Y(_645_) );
	NOR2X1 NOR2X1_45 ( .A(_525_), .B(_637_), .Y(_646_) );
	NAND2X1 NAND2X1_56 ( .A(_525_), .B(_637_), .Y(_647_) );
	OAI21X1 OAI21X1_237 ( .A(_645_), .B(_646_), .C(_647_), .Y(_648_) );
	OAI21X1 OAI21X1_238 ( .A(_633_), .B(_639_), .C(_648_), .Y(_649_) );
	XOR2X1 XOR2X1_6 ( .A(gen_nonce_synth_rand_10_), .B(_2__10_), .Y(_650_) );
	NAND2X1 NAND2X1_57 ( .A(_650_), .B(_649_), .Y(_651_) );
	INVX1 INVX1_198 ( .A(_649_), .Y(_652_) );
	INVX1 INVX1_199 ( .A(_650_), .Y(_653_) );
	NAND2X1 NAND2X1_58 ( .A(_653_), .B(_652_), .Y(_654_) );
	AOI21X1 AOI21X1_212 ( .A(_651_), .B(_654_), .C(comparador_valid_bF_buf0), .Y(_655_) );
	OAI21X1 OAI21X1_239 ( .A(_545__bF_buf4), .B(_2__10_), .C(_558__bF_buf2), .Y(_656_) );
	OAI22X1 OAI22X1_13 ( .A(_544_), .B(_644_), .C(_655_), .D(_656_), .Y(_517__10_) );
	INVX1 INVX1_200 ( .A(_2__11_), .Y(_657_) );
	OAI21X1 OAI21X1_240 ( .A(_526_), .B(_644_), .C(_651_), .Y(_658_) );
	XOR2X1 XOR2X1_7 ( .A(gen_nonce_synth_rand_11_), .B(_2__11_), .Y(_659_) );
	AND2X2 AND2X2_16 ( .A(_658_), .B(_659_), .Y(_660_) );
	OAI21X1 OAI21X1_241 ( .A(_658_), .B(_659_), .C(_545__bF_buf3), .Y(_661_) );
	OR2X2 OR2X2_11 ( .A(_660_), .B(_661_), .Y(_662_) );
	AOI21X1 AOI21X1_213 ( .A(comparador_valid_bF_buf5), .B(_2__11_), .C(_557_), .Y(_663_) );
	AOI22X1 AOI22X1_16 ( .A(_1__bF_buf5), .B(_657_), .C(_662_), .D(_663_), .Y(_517__11_) );
	NOR2X1 NOR2X1_46 ( .A(_2__12_), .B(_544_), .Y(_664_) );
	NOR2X1 NOR2X1_47 ( .A(_526_), .B(_644_), .Y(_665_) );
	NOR2X1 NOR2X1_48 ( .A(_527_), .B(_657_), .Y(_666_) );
	AOI21X1 AOI21X1_214 ( .A(_665_), .B(_659_), .C(_666_), .Y(_667_) );
	NAND2X1 NAND2X1_59 ( .A(_650_), .B(_659_), .Y(_668_) );
	OAI21X1 OAI21X1_242 ( .A(_668_), .B(_648_), .C(_667_), .Y(_669_) );
	NAND2X1 NAND2X1_60 ( .A(_632_), .B(_638_), .Y(_670_) );
	NOR2X1 NOR2X1_49 ( .A(_670_), .B(_668_), .Y(_671_) );
	AOI21X1 AOI21X1_215 ( .A(_671_), .B(_631_), .C(_669_), .Y(_672_) );
	XNOR2X1 XNOR2X1_8 ( .A(gen_nonce_synth_rand_12_), .B(_2__12_), .Y(_673_) );
	AOI21X1 AOI21X1_216 ( .A(_673_), .B(_672_), .C(comparador_valid_bF_buf4), .Y(_674_) );
	OAI21X1 OAI21X1_243 ( .A(_672_), .B(_673_), .C(_674_), .Y(_675_) );
	AOI21X1 AOI21X1_217 ( .A(comparador_valid_bF_buf3), .B(_2__12_), .C(_557_), .Y(_676_) );
	AOI21X1 AOI21X1_218 ( .A(_676_), .B(_675_), .C(_664_), .Y(_517__12_) );
	INVX1 INVX1_201 ( .A(_2__13_), .Y(_677_) );
	XNOR2X1 XNOR2X1_9 ( .A(gen_nonce_synth_rand_13_), .B(_2__13_), .Y(_678_) );
	NAND2X1 NAND2X1_61 ( .A(gen_nonce_synth_rand_12_), .B(_2__12_), .Y(_679_) );
	OAI21X1 OAI21X1_244 ( .A(_672_), .B(_673_), .C(_679_), .Y(_680_) );
	OAI21X1 OAI21X1_245 ( .A(_680_), .B(_678_), .C(_545__bF_buf2), .Y(_681_) );
	AOI21X1 AOI21X1_219 ( .A(_678_), .B(_680_), .C(_681_), .Y(_682_) );
	OAI21X1 OAI21X1_246 ( .A(_545__bF_buf1), .B(_2__13_), .C(_558__bF_buf1), .Y(_683_) );
	OAI22X1 OAI22X1_14 ( .A(_544_), .B(_677_), .C(_682_), .D(_683_), .Y(_517__13_) );
	INVX1 INVX1_202 ( .A(_2__14_), .Y(_684_) );
	XOR2X1 XOR2X1_8 ( .A(gen_nonce_synth_rand_12_), .B(_2__12_), .Y(_685_) );
	NAND2X1 NAND2X1_62 ( .A(gen_nonce_synth_rand_13_), .B(_2__13_), .Y(_686_) );
	NAND2X1 NAND2X1_63 ( .A(_529_), .B(_677_), .Y(_687_) );
	NAND3X1 NAND3X1_64 ( .A(_686_), .B(_687_), .C(_685_), .Y(_688_) );
	OAI21X1 OAI21X1_247 ( .A(_529_), .B(_677_), .C(_679_), .Y(_689_) );
	OAI21X1 OAI21X1_248 ( .A(gen_nonce_synth_rand_13_), .B(_2__13_), .C(_689_), .Y(_690_) );
	OAI21X1 OAI21X1_249 ( .A(_672_), .B(_688_), .C(_690_), .Y(_691_) );
	XOR2X1 XOR2X1_9 ( .A(gen_nonce_synth_rand_14_), .B(_2__14_), .Y(_692_) );
	AND2X2 AND2X2_17 ( .A(_691_), .B(_692_), .Y(_693_) );
	OAI21X1 OAI21X1_250 ( .A(_691_), .B(_692_), .C(_545__bF_buf0), .Y(_694_) );
	OR2X2 OR2X2_12 ( .A(_693_), .B(_694_), .Y(_695_) );
	AOI21X1 AOI21X1_220 ( .A(comparador_valid_bF_buf2), .B(_2__14_), .C(_557_), .Y(_696_) );
	AOI22X1 AOI22X1_17 ( .A(_1__bF_buf4), .B(_684_), .C(_695_), .D(_696_), .Y(_517__14_) );
	INVX1 INVX1_203 ( .A(_2__15_), .Y(_697_) );
	NOR2X1 NOR2X1_50 ( .A(_530_), .B(_684_), .Y(_698_) );
	NOR2X1 NOR2X1_51 ( .A(_698_), .B(_693_), .Y(_699_) );
	XNOR2X1 XNOR2X1_10 ( .A(gen_nonce_synth_rand_15_), .B(_2__15_), .Y(_700_) );
	AOI21X1 AOI21X1_221 ( .A(_700_), .B(_699_), .C(comparador_valid_bF_buf1), .Y(_701_) );
	OAI21X1 OAI21X1_251 ( .A(_699_), .B(_700_), .C(_701_), .Y(_702_) );
	AOI21X1 AOI21X1_222 ( .A(comparador_valid_bF_buf0), .B(_2__15_), .C(_557_), .Y(_703_) );
	AOI22X1 AOI22X1_18 ( .A(_1__bF_buf3), .B(_697_), .C(_702_), .D(_703_), .Y(_517__15_) );
	INVX1 INVX1_204 ( .A(_2__16_), .Y(_704_) );
	NOR2X1 NOR2X1_52 ( .A(_2__6_), .B(_523_), .Y(_705_) );
	NOR2X1 NOR2X1_53 ( .A(gen_nonce_synth_rand_6_), .B(_602_), .Y(_706_) );
	OAI21X1 OAI21X1_252 ( .A(_705_), .B(_706_), .C(_617_), .Y(_707_) );
	NOR2X1 NOR2X1_54 ( .A(_608_), .B(_707_), .Y(_708_) );
	OAI21X1 OAI21X1_253 ( .A(_589_), .B(_585_), .C(_708_), .Y(_709_) );
	XOR2X1 XOR2X1_10 ( .A(gen_nonce_synth_rand_15_), .B(_2__15_), .Y(_710_) );
	NAND2X1 NAND2X1_64 ( .A(_692_), .B(_710_), .Y(_711_) );
	NOR2X1 NOR2X1_55 ( .A(_711_), .B(_688_), .Y(_712_) );
	NAND2X1 NAND2X1_65 ( .A(_671_), .B(_712_), .Y(_713_) );
	AOI21X1 AOI21X1_223 ( .A(_630_), .B(_709_), .C(_713_), .Y(_714_) );
	NOR2X1 NOR2X1_56 ( .A(_531_), .B(_697_), .Y(_715_) );
	AOI21X1 AOI21X1_224 ( .A(_698_), .B(_710_), .C(_715_), .Y(_716_) );
	OAI21X1 OAI21X1_254 ( .A(_711_), .B(_690_), .C(_716_), .Y(_717_) );
	AOI21X1 AOI21X1_225 ( .A(_712_), .B(_669_), .C(_717_), .Y(_718_) );
	INVX1 INVX1_205 ( .A(_718_), .Y(_719_) );
	NOR2X1 NOR2X1_57 ( .A(_719_), .B(_714_), .Y(_720_) );
	NAND2X1 NAND2X1_66 ( .A(gen_nonce_synth_rand_16_), .B(_2__16_), .Y(_721_) );
	NAND2X1 NAND2X1_67 ( .A(_532_), .B(_704_), .Y(_722_) );
	NAND2X1 NAND2X1_68 ( .A(_721_), .B(_722_), .Y(_723_) );
	AOI21X1 AOI21X1_226 ( .A(_723_), .B(_720_), .C(comparador_valid_bF_buf5), .Y(_724_) );
	OAI21X1 OAI21X1_255 ( .A(_720_), .B(_723_), .C(_724_), .Y(_725_) );
	AOI21X1 AOI21X1_227 ( .A(comparador_valid_bF_buf4), .B(_2__16_), .C(_557_), .Y(_726_) );
	AOI22X1 AOI22X1_19 ( .A(_1__bF_buf2), .B(_704_), .C(_725_), .D(_726_), .Y(_517__16_) );
	INVX1 INVX1_206 ( .A(_2__17_), .Y(_727_) );
	OAI21X1 OAI21X1_256 ( .A(_720_), .B(_723_), .C(_721_), .Y(_728_) );
	NOR2X1 NOR2X1_58 ( .A(_533_), .B(_727_), .Y(_729_) );
	NOR2X1 NOR2X1_59 ( .A(gen_nonce_synth_rand_17_), .B(_2__17_), .Y(_730_) );
	OR2X2 OR2X2_13 ( .A(_729_), .B(_730_), .Y(_731_) );
	OAI21X1 OAI21X1_257 ( .A(_728_), .B(_731_), .C(_545__bF_buf4), .Y(_732_) );
	AOI21X1 AOI21X1_228 ( .A(_728_), .B(_731_), .C(_732_), .Y(_733_) );
	OAI21X1 OAI21X1_258 ( .A(_545__bF_buf3), .B(_2__17_), .C(_558__bF_buf0), .Y(_734_) );
	OAI22X1 OAI22X1_15 ( .A(_544_), .B(_727_), .C(_733_), .D(_734_), .Y(_517__17_) );
	INVX1 INVX1_207 ( .A(_2__18_), .Y(_735_) );
	OAI21X1 OAI21X1_259 ( .A(_533_), .B(_727_), .C(_721_), .Y(_736_) );
	OAI21X1 OAI21X1_260 ( .A(gen_nonce_synth_rand_17_), .B(_2__17_), .C(_736_), .Y(_737_) );
	NOR2X1 NOR2X1_60 ( .A(_723_), .B(_731_), .Y(_738_) );
	INVX1 INVX1_208 ( .A(_738_), .Y(_739_) );
	OAI21X1 OAI21X1_261 ( .A(_720_), .B(_739_), .C(_737_), .Y(_740_) );
	NAND2X1 NAND2X1_69 ( .A(gen_nonce_synth_rand_18_), .B(_2__18_), .Y(_741_) );
	NAND2X1 NAND2X1_70 ( .A(_534_), .B(_735_), .Y(_742_) );
	AND2X2 AND2X2_18 ( .A(_742_), .B(_741_), .Y(_743_) );
	OR2X2 OR2X2_14 ( .A(_740_), .B(_743_), .Y(_744_) );
	NAND2X1 NAND2X1_71 ( .A(_743_), .B(_740_), .Y(_745_) );
	AOI21X1 AOI21X1_229 ( .A(_745_), .B(_744_), .C(comparador_valid_bF_buf3), .Y(_746_) );
	OAI21X1 OAI21X1_262 ( .A(_545__bF_buf2), .B(_2__18_), .C(_558__bF_buf3), .Y(_747_) );
	OAI22X1 OAI22X1_16 ( .A(_544_), .B(_735_), .C(_746_), .D(_747_), .Y(_517__18_) );
	INVX1 INVX1_209 ( .A(_2__19_), .Y(_748_) );
	AND2X2 AND2X2_19 ( .A(_745_), .B(_741_), .Y(_749_) );
	NAND2X1 NAND2X1_72 ( .A(gen_nonce_synth_rand_19_), .B(_2__19_), .Y(_750_) );
	NAND2X1 NAND2X1_73 ( .A(_535_), .B(_748_), .Y(_751_) );
	NAND2X1 NAND2X1_74 ( .A(_750_), .B(_751_), .Y(_752_) );
	AOI21X1 AOI21X1_230 ( .A(_752_), .B(_749_), .C(comparador_valid_bF_buf2), .Y(_753_) );
	OAI21X1 OAI21X1_263 ( .A(_749_), .B(_752_), .C(_753_), .Y(_754_) );
	AOI21X1 AOI21X1_231 ( .A(comparador_valid_bF_buf1), .B(_2__19_), .C(_557_), .Y(_755_) );
	AOI22X1 AOI22X1_20 ( .A(_1__bF_buf1), .B(_748_), .C(_754_), .D(_755_), .Y(_517__19_) );
	INVX1 INVX1_210 ( .A(_2__20_), .Y(_756_) );
	INVX1 INVX1_211 ( .A(_737_), .Y(_757_) );
	NAND2X1 NAND2X1_75 ( .A(_741_), .B(_742_), .Y(_758_) );
	NOR2X1 NOR2X1_61 ( .A(_758_), .B(_752_), .Y(_759_) );
	OAI21X1 OAI21X1_264 ( .A(_752_), .B(_741_), .C(_750_), .Y(_760_) );
	AOI21X1 AOI21X1_232 ( .A(_759_), .B(_757_), .C(_760_), .Y(_761_) );
	NAND2X1 NAND2X1_76 ( .A(_759_), .B(_738_), .Y(_762_) );
	OAI21X1 OAI21X1_265 ( .A(_720_), .B(_762_), .C(_761_), .Y(_763_) );
	XOR2X1 XOR2X1_11 ( .A(gen_nonce_synth_rand_20_), .B(_2__20_), .Y(_764_) );
	NAND2X1 NAND2X1_77 ( .A(_764_), .B(_763_), .Y(_765_) );
	OR2X2 OR2X2_15 ( .A(_763_), .B(_764_), .Y(_766_) );
	AOI21X1 AOI21X1_233 ( .A(_765_), .B(_766_), .C(comparador_valid_bF_buf0), .Y(_767_) );
	OAI21X1 OAI21X1_266 ( .A(_545__bF_buf1), .B(_2__20_), .C(_558__bF_buf2), .Y(_768_) );
	OAI22X1 OAI22X1_17 ( .A(_544_), .B(_756_), .C(_767_), .D(_768_), .Y(_517__20_) );
	INVX1 INVX1_212 ( .A(_2__21_), .Y(_769_) );
	OAI21X1 OAI21X1_267 ( .A(_536_), .B(_756_), .C(_765_), .Y(_770_) );
	NOR2X1 NOR2X1_62 ( .A(_537_), .B(_769_), .Y(_771_) );
	NOR2X1 NOR2X1_63 ( .A(gen_nonce_synth_rand_21_), .B(_2__21_), .Y(_772_) );
	NOR2X1 NOR2X1_64 ( .A(_772_), .B(_771_), .Y(_773_) );
	NAND2X1 NAND2X1_78 ( .A(_773_), .B(_770_), .Y(_774_) );
	OR2X2 OR2X2_16 ( .A(_770_), .B(_773_), .Y(_775_) );
	NAND3X1 NAND3X1_65 ( .A(_545__bF_buf0), .B(_774_), .C(_775_), .Y(_776_) );
	AOI21X1 AOI21X1_234 ( .A(comparador_valid_bF_buf5), .B(_2__21_), .C(_557_), .Y(_777_) );
	AOI22X1 AOI22X1_21 ( .A(_1__bF_buf0), .B(_769_), .C(_776_), .D(_777_), .Y(_517__21_) );
	NAND2X1 NAND2X1_79 ( .A(_1__bF_buf5), .B(_2__22_), .Y(_778_) );
	NAND2X1 NAND2X1_80 ( .A(gen_nonce_synth_rand_22_), .B(_2__22_), .Y(_779_) );
	INVX1 INVX1_213 ( .A(_779_), .Y(_780_) );
	NOR2X1 NOR2X1_65 ( .A(gen_nonce_synth_rand_22_), .B(_2__22_), .Y(_781_) );
	OR2X2 OR2X2_17 ( .A(_780_), .B(_781_), .Y(_782_) );
	AND2X2 AND2X2_20 ( .A(_773_), .B(_764_), .Y(_783_) );
	NAND2X1 NAND2X1_81 ( .A(_783_), .B(_763_), .Y(_784_) );
	NAND2X1 NAND2X1_82 ( .A(gen_nonce_synth_rand_20_), .B(_2__20_), .Y(_785_) );
	INVX1 INVX1_214 ( .A(_771_), .Y(_786_) );
	OAI21X1 OAI21X1_268 ( .A(_772_), .B(_785_), .C(_786_), .Y(_787_) );
	INVX1 INVX1_215 ( .A(_787_), .Y(_788_) );
	NAND3X1 NAND3X1_66 ( .A(_782_), .B(_788_), .C(_784_), .Y(_789_) );
	INVX1 INVX1_216 ( .A(_782_), .Y(_790_) );
	AND2X2 AND2X2_21 ( .A(_763_), .B(_783_), .Y(_791_) );
	OAI21X1 OAI21X1_269 ( .A(_791_), .B(_787_), .C(_790_), .Y(_792_) );
	AOI21X1 AOI21X1_235 ( .A(_789_), .B(_792_), .C(comparador_valid_bF_buf4), .Y(_793_) );
	OAI21X1 OAI21X1_270 ( .A(_545__bF_buf4), .B(_2__22_), .C(_558__bF_buf1), .Y(_794_) );
	OAI21X1 OAI21X1_271 ( .A(_793_), .B(_794_), .C(_778_), .Y(_517__22_) );
	INVX1 INVX1_217 ( .A(_2__23_), .Y(_795_) );
	AOI21X1 AOI21X1_236 ( .A(_788_), .B(_784_), .C(_782_), .Y(_796_) );
	NOR2X1 NOR2X1_66 ( .A(_539_), .B(_795_), .Y(_797_) );
	NOR2X1 NOR2X1_67 ( .A(gen_nonce_synth_rand_23_), .B(_2__23_), .Y(_798_) );
	OR2X2 OR2X2_18 ( .A(_797_), .B(_798_), .Y(_799_) );
	INVX1 INVX1_218 ( .A(_799_), .Y(_800_) );
	OAI21X1 OAI21X1_272 ( .A(_796_), .B(_780_), .C(_800_), .Y(_801_) );
	NAND3X1 NAND3X1_67 ( .A(_779_), .B(_799_), .C(_792_), .Y(_802_) );
	NAND3X1 NAND3X1_68 ( .A(_545__bF_buf3), .B(_801_), .C(_802_), .Y(_803_) );
	AOI21X1 AOI21X1_237 ( .A(comparador_valid_bF_buf3), .B(_2__23_), .C(_557_), .Y(_804_) );
	AOI22X1 AOI22X1_22 ( .A(_1__bF_buf4), .B(_795_), .C(_803_), .D(_804_), .Y(_517__23_) );
	INVX1 INVX1_219 ( .A(_2__24_), .Y(_805_) );
	NAND2X1 NAND2X1_83 ( .A(gen_nonce_synth_rand_8_), .B(_623_), .Y(_806_) );
	NAND2X1 NAND2X1_84 ( .A(_2__8_), .B(_524_), .Y(_807_) );
	NAND2X1 NAND2X1_85 ( .A(gen_nonce_synth_rand_9_), .B(_637_), .Y(_808_) );
	NAND2X1 NAND2X1_86 ( .A(_2__9_), .B(_525_), .Y(_809_) );
	AOI22X1 AOI22X1_23 ( .A(_806_), .B(_807_), .C(_808_), .D(_809_), .Y(_810_) );
	NAND3X1 NAND3X1_69 ( .A(_650_), .B(_659_), .C(_810_), .Y(_811_) );
	NOR3X1 NOR3X1_2 ( .A(_688_), .B(_711_), .C(_811_), .Y(_812_) );
	NAND2X1 NAND2X1_87 ( .A(_631_), .B(_812_), .Y(_813_) );
	NOR2X1 NOR2X1_68 ( .A(_782_), .B(_799_), .Y(_814_) );
	NAND2X1 NAND2X1_88 ( .A(_783_), .B(_814_), .Y(_815_) );
	OR2X2 OR2X2_19 ( .A(_762_), .B(_815_), .Y(_816_) );
	AOI21X1 AOI21X1_238 ( .A(_718_), .B(_813_), .C(_816_), .Y(_817_) );
	NOR2X1 NOR2X1_69 ( .A(_761_), .B(_815_), .Y(_818_) );
	AOI21X1 AOI21X1_239 ( .A(_780_), .B(_800_), .C(_797_), .Y(_819_) );
	NAND2X1 NAND2X1_89 ( .A(_787_), .B(_814_), .Y(_820_) );
	NAND2X1 NAND2X1_90 ( .A(_819_), .B(_820_), .Y(_821_) );
	OR2X2 OR2X2_20 ( .A(_818_), .B(_821_), .Y(_822_) );
	NOR2X1 NOR2X1_70 ( .A(_540_), .B(_805_), .Y(_823_) );
	INVX1 INVX1_220 ( .A(_823_), .Y(_824_) );
	NAND2X1 NAND2X1_91 ( .A(_540_), .B(_805_), .Y(_825_) );
	NAND2X1 NAND2X1_92 ( .A(_825_), .B(_824_), .Y(_826_) );
	INVX1 INVX1_221 ( .A(_826_), .Y(_827_) );
	OAI21X1 OAI21X1_273 ( .A(_817_), .B(_822_), .C(_827_), .Y(_828_) );
	NOR2X1 NOR2X1_71 ( .A(_822_), .B(_817_), .Y(_829_) );
	NAND2X1 NAND2X1_93 ( .A(_826_), .B(_829_), .Y(_830_) );
	AOI21X1 AOI21X1_240 ( .A(_828_), .B(_830_), .C(comparador_valid_bF_buf2), .Y(_831_) );
	OAI21X1 OAI21X1_274 ( .A(_545__bF_buf2), .B(_2__24_), .C(_558__bF_buf0), .Y(_832_) );
	OAI22X1 OAI22X1_18 ( .A(_544_), .B(_805_), .C(_831_), .D(_832_), .Y(_517__24_) );
	NAND2X1 NAND2X1_94 ( .A(_1__bF_buf3), .B(_2__25_), .Y(_833_) );
	NAND2X1 NAND2X1_95 ( .A(gen_nonce_synth_rand_25_), .B(_2__25_), .Y(_834_) );
	INVX1 INVX1_222 ( .A(_834_), .Y(_835_) );
	NOR2X1 NOR2X1_72 ( .A(gen_nonce_synth_rand_25_), .B(_2__25_), .Y(_836_) );
	NOR2X1 NOR2X1_73 ( .A(_836_), .B(_835_), .Y(_837_) );
	OAI21X1 OAI21X1_275 ( .A(_540_), .B(_805_), .C(_828_), .Y(_838_) );
	OR2X2 OR2X2_21 ( .A(_838_), .B(_837_), .Y(_839_) );
	INVX1 INVX1_223 ( .A(_837_), .Y(_840_) );
	NOR2X1 NOR2X1_74 ( .A(_826_), .B(_840_), .Y(_841_) );
	OAI21X1 OAI21X1_276 ( .A(_817_), .B(_822_), .C(_841_), .Y(_842_) );
	OAI21X1 OAI21X1_277 ( .A(_824_), .B(_840_), .C(_842_), .Y(_843_) );
	INVX1 INVX1_224 ( .A(_843_), .Y(_844_) );
	AOI21X1 AOI21X1_241 ( .A(_844_), .B(_839_), .C(comparador_valid_bF_buf1), .Y(_845_) );
	OAI21X1 OAI21X1_278 ( .A(_545__bF_buf1), .B(_2__25_), .C(_558__bF_buf3), .Y(_846_) );
	OAI21X1 OAI21X1_279 ( .A(_845_), .B(_846_), .C(_833_), .Y(_517__25_) );
	NAND2X1 NAND2X1_96 ( .A(_1__bF_buf2), .B(_2__26_), .Y(_847_) );
	OAI21X1 OAI21X1_280 ( .A(_824_), .B(_836_), .C(_834_), .Y(_848_) );
	INVX1 INVX1_225 ( .A(_848_), .Y(_849_) );
	XNOR2X1 XNOR2X1_11 ( .A(gen_nonce_synth_rand_26_), .B(_2__26_), .Y(_850_) );
	NAND3X1 NAND3X1_70 ( .A(_849_), .B(_850_), .C(_842_), .Y(_851_) );
	AOI21X1 AOI21X1_242 ( .A(_849_), .B(_842_), .C(_850_), .Y(_852_) );
	INVX1 INVX1_226 ( .A(_852_), .Y(_853_) );
	AOI21X1 AOI21X1_243 ( .A(_851_), .B(_853_), .C(comparador_valid_bF_buf0), .Y(_854_) );
	OAI21X1 OAI21X1_281 ( .A(_545__bF_buf0), .B(_2__26_), .C(_558__bF_buf2), .Y(_855_) );
	OAI21X1 OAI21X1_282 ( .A(_854_), .B(_855_), .C(_847_), .Y(_517__26_) );
	NAND2X1 NAND2X1_97 ( .A(gen_nonce_synth_rand_26_), .B(_2__26_), .Y(_856_) );
	INVX1 INVX1_227 ( .A(_856_), .Y(_857_) );
	NAND2X1 NAND2X1_98 ( .A(gen_nonce_synth_rand_27_), .B(_2__27_), .Y(_858_) );
	INVX1 INVX1_228 ( .A(_858_), .Y(_859_) );
	NOR2X1 NOR2X1_75 ( .A(gen_nonce_synth_rand_27_), .B(_2__27_), .Y(_860_) );
	NOR2X1 NOR2X1_76 ( .A(_860_), .B(_859_), .Y(_861_) );
	OAI21X1 OAI21X1_283 ( .A(_852_), .B(_857_), .C(_861_), .Y(_862_) );
	NOR2X1 NOR2X1_77 ( .A(_857_), .B(_852_), .Y(_863_) );
	OAI21X1 OAI21X1_284 ( .A(_859_), .B(_860_), .C(_863_), .Y(_864_) );
	AOI21X1 AOI21X1_244 ( .A(_862_), .B(_864_), .C(comparador_valid_bF_buf5), .Y(_865_) );
	OAI21X1 OAI21X1_285 ( .A(_545__bF_buf4), .B(_2__27_), .C(_558__bF_buf1), .Y(_866_) );
	NAND2X1 NAND2X1_99 ( .A(_1__bF_buf1), .B(_2__27_), .Y(_867_) );
	OAI21X1 OAI21X1_286 ( .A(_865_), .B(_866_), .C(_867_), .Y(_517__27_) );
	INVX1 INVX1_229 ( .A(_2__28_), .Y(_868_) );
	INVX1 INVX1_230 ( .A(_850_), .Y(_869_) );
	NAND2X1 NAND2X1_100 ( .A(_861_), .B(_869_), .Y(_870_) );
	INVX1 INVX1_231 ( .A(_870_), .Y(_871_) );
	NAND2X1 NAND2X1_101 ( .A(_871_), .B(_841_), .Y(_872_) );
	OAI21X1 OAI21X1_287 ( .A(_860_), .B(_856_), .C(_858_), .Y(_873_) );
	INVX1 INVX1_232 ( .A(_873_), .Y(_874_) );
	OAI21X1 OAI21X1_288 ( .A(_849_), .B(_870_), .C(_874_), .Y(_875_) );
	INVX1 INVX1_233 ( .A(_875_), .Y(_876_) );
	OAI21X1 OAI21X1_289 ( .A(_829_), .B(_872_), .C(_876_), .Y(_877_) );
	NOR2X1 NOR2X1_78 ( .A(_542_), .B(_868_), .Y(_878_) );
	INVX1 INVX1_234 ( .A(_878_), .Y(_879_) );
	NAND2X1 NAND2X1_102 ( .A(_542_), .B(_868_), .Y(_880_) );
	AND2X2 AND2X2_22 ( .A(_879_), .B(_880_), .Y(_881_) );
	NOR2X1 NOR2X1_79 ( .A(_881_), .B(_877_), .Y(_882_) );
	NOR2X1 NOR2X1_80 ( .A(_762_), .B(_815_), .Y(_883_) );
	OAI21X1 OAI21X1_290 ( .A(_714_), .B(_719_), .C(_883_), .Y(_884_) );
	NOR2X1 NOR2X1_81 ( .A(_821_), .B(_818_), .Y(_885_) );
	AOI21X1 AOI21X1_245 ( .A(_885_), .B(_884_), .C(_872_), .Y(_886_) );
	OAI21X1 OAI21X1_291 ( .A(_886_), .B(_875_), .C(_881_), .Y(_887_) );
	INVX1 INVX1_235 ( .A(_887_), .Y(_888_) );
	OAI21X1 OAI21X1_292 ( .A(_882_), .B(_888_), .C(_545__bF_buf3), .Y(_889_) );
	OAI21X1 OAI21X1_293 ( .A(_545__bF_buf2), .B(_2__28_), .C(_889_), .Y(_890_) );
	OAI22X1 OAI22X1_19 ( .A(_544_), .B(_868_), .C(_890_), .D(_557_), .Y(_517__28_) );
	INVX1 INVX1_236 ( .A(_2__29_), .Y(_891_) );
	OAI21X1 OAI21X1_294 ( .A(_542_), .B(_868_), .C(_887_), .Y(_892_) );
	NOR2X1 NOR2X1_82 ( .A(_543_), .B(_891_), .Y(_893_) );
	NOR2X1 NOR2X1_83 ( .A(gen_nonce_synth_rand_29_), .B(_2__29_), .Y(_894_) );
	NOR2X1 NOR2X1_84 ( .A(_894_), .B(_893_), .Y(_895_) );
	INVX1 INVX1_237 ( .A(_895_), .Y(_896_) );
	OAI21X1 OAI21X1_295 ( .A(_892_), .B(_896_), .C(_545__bF_buf1), .Y(_897_) );
	AOI21X1 AOI21X1_246 ( .A(_892_), .B(_896_), .C(_897_), .Y(_898_) );
	OAI21X1 OAI21X1_296 ( .A(_545__bF_buf0), .B(_2__29_), .C(_558__bF_buf0), .Y(_899_) );
	OAI22X1 OAI22X1_20 ( .A(_544_), .B(_891_), .C(_898_), .D(_899_), .Y(_517__29_) );
	NAND2X1 NAND2X1_103 ( .A(_1__bF_buf0), .B(_2__30_), .Y(_900_) );
	INVX1 INVX1_238 ( .A(_872_), .Y(_901_) );
	OAI21X1 OAI21X1_297 ( .A(_817_), .B(_822_), .C(_901_), .Y(_902_) );
	INVX1 INVX1_239 ( .A(_881_), .Y(_903_) );
	NOR2X1 NOR2X1_85 ( .A(_896_), .B(_903_), .Y(_904_) );
	INVX1 INVX1_240 ( .A(_904_), .Y(_905_) );
	AOI21X1 AOI21X1_247 ( .A(_876_), .B(_902_), .C(_905_), .Y(_906_) );
	AOI21X1 AOI21X1_248 ( .A(_878_), .B(_895_), .C(_893_), .Y(_907_) );
	INVX1 INVX1_241 ( .A(_907_), .Y(_908_) );
	NAND2X1 NAND2X1_104 ( .A(gen_nonce_synth_rand_30_), .B(_2__30_), .Y(_909_) );
	INVX1 INVX1_242 ( .A(_909_), .Y(_910_) );
	NOR2X1 NOR2X1_86 ( .A(gen_nonce_synth_rand_30_), .B(_2__30_), .Y(_911_) );
	NOR2X1 NOR2X1_87 ( .A(_911_), .B(_910_), .Y(_912_) );
	OAI21X1 OAI21X1_298 ( .A(_906_), .B(_908_), .C(_912_), .Y(_913_) );
	OAI21X1 OAI21X1_299 ( .A(_886_), .B(_875_), .C(_904_), .Y(_914_) );
	INVX1 INVX1_243 ( .A(_912_), .Y(_915_) );
	NAND3X1 NAND3X1_71 ( .A(_907_), .B(_915_), .C(_914_), .Y(_916_) );
	AOI21X1 AOI21X1_249 ( .A(_916_), .B(_913_), .C(comparador_valid_bF_buf4), .Y(_917_) );
	OAI21X1 OAI21X1_300 ( .A(_545__bF_buf4), .B(_2__30_), .C(_558__bF_buf3), .Y(_918_) );
	OAI21X1 OAI21X1_301 ( .A(_917_), .B(_918_), .C(_900_), .Y(_517__30_) );
	AOI21X1 AOI21X1_250 ( .A(_907_), .B(_914_), .C(_915_), .Y(_919_) );
	XNOR2X1 XNOR2X1_12 ( .A(gen_nonce_synth_rand_31_), .B(_2__31_), .Y(_920_) );
	INVX1 INVX1_244 ( .A(_920_), .Y(_921_) );
	OAI21X1 OAI21X1_302 ( .A(_919_), .B(_910_), .C(_921_), .Y(_922_) );
	NAND3X1 NAND3X1_72 ( .A(_909_), .B(_920_), .C(_913_), .Y(_923_) );
	NAND3X1 NAND3X1_73 ( .A(_545__bF_buf3), .B(_923_), .C(_922_), .Y(_924_) );
	AOI21X1 AOI21X1_251 ( .A(comparador_valid_bF_buf3), .B(_2__31_), .C(_557_), .Y(_925_) );
	NOR2X1 NOR2X1_88 ( .A(_2__31_), .B(_544_), .Y(_926_) );
	AOI21X1 AOI21X1_252 ( .A(_925_), .B(_924_), .C(_926_), .Y(_517__31_) );
	DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf31), .D(_517__0_), .Q(_2__0_) );
	DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf30), .D(_517__1_), .Q(_2__1_) );
	DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf29), .D(_517__2_), .Q(_2__2_) );
	DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf28), .D(_517__3_), .Q(_2__3_) );
	DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf27), .D(_517__4_), .Q(_2__4_) );
	DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf26), .D(_517__5_), .Q(_2__5_) );
	DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf25), .D(_517__6_), .Q(_2__6_) );
	DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf24), .D(_517__7_), .Q(_2__7_) );
	DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf23), .D(_517__8_), .Q(_2__8_) );
	DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf22), .D(_517__9_), .Q(_2__9_) );
	DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf21), .D(_517__10_), .Q(_2__10_) );
	DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf20), .D(_517__11_), .Q(_2__11_) );
	DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf19), .D(_517__12_), .Q(_2__12_) );
	DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf18), .D(_517__13_), .Q(_2__13_) );
	DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf17), .D(_517__14_), .Q(_2__14_) );
	DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf16), .D(_517__15_), .Q(_2__15_) );
	DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf15), .D(_517__16_), .Q(_2__16_) );
	DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf14), .D(_517__17_), .Q(_2__17_) );
	DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf13), .D(_517__18_), .Q(_2__18_) );
	DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf12), .D(_517__19_), .Q(_2__19_) );
	DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf11), .D(_517__20_), .Q(_2__20_) );
	DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf10), .D(_517__21_), .Q(_2__21_) );
	DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf9), .D(_517__22_), .Q(_2__22_) );
	DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf8), .D(_517__23_), .Q(_2__23_) );
	DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf7), .D(_517__24_), .Q(_2__24_) );
	DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf6), .D(_517__25_), .Q(_2__25_) );
	DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf5), .D(_517__26_), .Q(_2__26_) );
	DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf4), .D(_517__27_), .Q(_2__27_) );
	DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf3), .D(_517__28_), .Q(_2__28_) );
	DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf2), .D(_517__29_), .Q(_2__29_) );
	DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf1), .D(_517__30_), .Q(_2__30_) );
	DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf0), .D(_517__31_), .Q(_2__31_) );
	DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf76), .D(_518__0_), .Q(gen_nonce_synth_rand_0_) );
	DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf75), .D(_518__1_), .Q(gen_nonce_synth_rand_1_) );
	DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf74), .D(_518__2_), .Q(gen_nonce_synth_rand_2_) );
	DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf73), .D(_518__3_), .Q(gen_nonce_synth_rand_3_) );
	DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf72), .D(_518__4_), .Q(gen_nonce_synth_rand_4_) );
	DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf71), .D(_518__5_), .Q(gen_nonce_synth_rand_5_) );
	DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf70), .D(_518__6_), .Q(gen_nonce_synth_rand_6_) );
	DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf69), .D(_518__7_), .Q(gen_nonce_synth_rand_7_) );
	DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf68), .D(_518__8_), .Q(gen_nonce_synth_rand_8_) );
	DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf67), .D(_518__9_), .Q(gen_nonce_synth_rand_9_) );
	DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf66), .D(_518__10_), .Q(gen_nonce_synth_rand_10_) );
	DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf65), .D(_518__11_), .Q(gen_nonce_synth_rand_11_) );
	DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf64), .D(_518__12_), .Q(gen_nonce_synth_rand_12_) );
	DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf63), .D(_518__13_), .Q(gen_nonce_synth_rand_13_) );
	DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf62), .D(_518__14_), .Q(gen_nonce_synth_rand_14_) );
	DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf61), .D(_518__15_), .Q(gen_nonce_synth_rand_15_) );
	DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf60), .D(_518__16_), .Q(gen_nonce_synth_rand_16_) );
	DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf59), .D(_518__17_), .Q(gen_nonce_synth_rand_17_) );
	DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf58), .D(_518__18_), .Q(gen_nonce_synth_rand_18_) );
	DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf57), .D(_518__19_), .Q(gen_nonce_synth_rand_19_) );
	DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf56), .D(_518__20_), .Q(gen_nonce_synth_rand_20_) );
	DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf55), .D(_518__21_), .Q(gen_nonce_synth_rand_21_) );
	DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf54), .D(_518__22_), .Q(gen_nonce_synth_rand_22_) );
	DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf53), .D(_518__23_), .Q(gen_nonce_synth_rand_23_) );
	DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf52), .D(_518__24_), .Q(gen_nonce_synth_rand_24_) );
	DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf51), .D(_518__25_), .Q(gen_nonce_synth_rand_25_) );
	DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf50), .D(_518__26_), .Q(gen_nonce_synth_rand_26_) );
	DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf49), .D(_518__27_), .Q(gen_nonce_synth_rand_27_) );
	DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf48), .D(_518__28_), .Q(gen_nonce_synth_rand_28_) );
	DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf47), .D(_518__29_), .Q(gen_nonce_synth_rand_29_) );
	DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf46), .D(_518__30_), .Q(gen_nonce_synth_rand_30_) );
	DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf45), .D(_518__31_), .Q(gen_nonce_synth_rand_31_) );
	INVX1 INVX1_245 ( .A(micro_hash_synth_W_27__0_), .Y(_2461_) );
	INVX1 INVX1_246 ( .A(concatenador_count_0_bF_buf10), .Y(_2462_) );
	INVX4 INVX4_3 ( .A(concatenador_count_1_bF_buf5), .Y(_2463_) );
	NOR2X1 NOR2X1_89 ( .A(concatenador_count_3_), .B(concatenador_count_2_), .Y(_2464_) );
	INVX1 INVX1_247 ( .A(_2464_), .Y(_2465_) );
	NOR2X1 NOR2X1_90 ( .A(concatenador_count_4_), .B(_2465_), .Y(_2466_) );
	OAI21X1 OAI21X1_303 ( .A(_2462_), .B(_2463_), .C(_2466_), .Y(_2467_) );
	NOR2X1 NOR2X1_91 ( .A(concatenador_count_5_), .B(_2467_), .Y(_2468_) );
	INVX1 INVX1_248 ( .A(_2468_), .Y(_2469_) );
	NOR2X1 NOR2X1_92 ( .A(concatenador_count_0_bF_buf9), .B(concatenador_count_1_bF_buf4), .Y(_2470_) );
	OAI21X1 OAI21X1_304 ( .A(_2469_), .B(_2470__bF_buf3), .C(reset_L_bF_buf5), .Y(_2471_) );
	NOR2X1 NOR2X1_93 ( .A(_2470__bF_buf2), .B(_2469_), .Y(_2472_) );
	NAND2X1 NAND2X1_105 ( .A(reset_L_bF_buf4), .B(_2472_), .Y(_2473_) );
	INVX1 INVX1_249 ( .A(micro_hash_synth_W_13__0_), .Y(_2474_) );
	INVX1 INVX1_250 ( .A(micro_hash_synth_W_24__0_), .Y(_2475_) );
	OAI21X1 OAI21X1_305 ( .A(_2474_), .B(micro_hash_synth_W_18__0_), .C(_2475_), .Y(_2476_) );
	AOI21X1 AOI21X1_253 ( .A(_2474_), .B(micro_hash_synth_W_18__0_), .C(_2476_), .Y(_2477_) );
	OAI22X1 OAI22X1_21 ( .A(_2461_), .B(_2471__bF_buf13), .C(_2473__bF_buf15), .D(_2477_), .Y(_1109_) );
	INVX1 INVX1_251 ( .A(micro_hash_synth_W_27__1_), .Y(_2478_) );
	INVX1 INVX1_252 ( .A(micro_hash_synth_W_13__1_), .Y(_2479_) );
	INVX1 INVX1_253 ( .A(micro_hash_synth_W_24__1_), .Y(_2480_) );
	OAI21X1 OAI21X1_306 ( .A(_2479_), .B(micro_hash_synth_W_18__1_), .C(_2480_), .Y(_2481_) );
	AOI21X1 AOI21X1_254 ( .A(_2479_), .B(micro_hash_synth_W_18__1_), .C(_2481_), .Y(_2482_) );
	OAI22X1 OAI22X1_22 ( .A(_2478_), .B(_2471__bF_buf12), .C(_2473__bF_buf14), .D(_2482_), .Y(_1110_) );
	INVX1 INVX1_254 ( .A(micro_hash_synth_W_27__2_), .Y(_2483_) );
	INVX1 INVX1_255 ( .A(micro_hash_synth_W_13__2_), .Y(_2484_) );
	INVX1 INVX1_256 ( .A(micro_hash_synth_W_24__2_), .Y(_2485_) );
	OAI21X1 OAI21X1_307 ( .A(_2484_), .B(micro_hash_synth_W_18__2_), .C(_2485_), .Y(_2486_) );
	AOI21X1 AOI21X1_255 ( .A(_2484_), .B(micro_hash_synth_W_18__2_), .C(_2486_), .Y(_2487_) );
	OAI22X1 OAI22X1_23 ( .A(_2483_), .B(_2471__bF_buf11), .C(_2473__bF_buf13), .D(_2487_), .Y(_1111_) );
	INVX1 INVX1_257 ( .A(micro_hash_synth_W_27__3_), .Y(_2488_) );
	INVX1 INVX1_258 ( .A(micro_hash_synth_W_13__3_), .Y(_2489_) );
	INVX1 INVX1_259 ( .A(micro_hash_synth_W_24__3_), .Y(_2490_) );
	OAI21X1 OAI21X1_308 ( .A(_2489_), .B(micro_hash_synth_W_18__3_), .C(_2490_), .Y(_2491_) );
	AOI21X1 AOI21X1_256 ( .A(_2489_), .B(micro_hash_synth_W_18__3_), .C(_2491_), .Y(_2492_) );
	OAI22X1 OAI22X1_24 ( .A(_2488_), .B(_2471__bF_buf10), .C(_2473__bF_buf12), .D(_2492_), .Y(_1112_) );
	INVX1 INVX1_260 ( .A(micro_hash_synth_W_27__4_), .Y(_2493_) );
	INVX1 INVX1_261 ( .A(micro_hash_synth_W_13__4_), .Y(_2494_) );
	INVX1 INVX1_262 ( .A(micro_hash_synth_W_24__4_), .Y(_2495_) );
	OAI21X1 OAI21X1_309 ( .A(_2494_), .B(micro_hash_synth_W_18__4_), .C(_2495_), .Y(_2496_) );
	AOI21X1 AOI21X1_257 ( .A(_2494_), .B(micro_hash_synth_W_18__4_), .C(_2496_), .Y(_2497_) );
	OAI22X1 OAI22X1_25 ( .A(_2493_), .B(_2471__bF_buf9), .C(_2473__bF_buf11), .D(_2497_), .Y(_1113_) );
	INVX1 INVX1_263 ( .A(micro_hash_synth_W_27__5_), .Y(_2498_) );
	INVX1 INVX1_264 ( .A(micro_hash_synth_W_13__5_), .Y(_2499_) );
	INVX1 INVX1_265 ( .A(micro_hash_synth_W_24__5_), .Y(_2500_) );
	OAI21X1 OAI21X1_310 ( .A(_2499_), .B(micro_hash_synth_W_18__5_), .C(_2500_), .Y(_2501_) );
	AOI21X1 AOI21X1_258 ( .A(_2499_), .B(micro_hash_synth_W_18__5_), .C(_2501_), .Y(_2502_) );
	OAI22X1 OAI22X1_26 ( .A(_2498_), .B(_2471__bF_buf8), .C(_2473__bF_buf10), .D(_2502_), .Y(_1114_) );
	INVX1 INVX1_266 ( .A(micro_hash_synth_W_27__6_), .Y(_2503_) );
	INVX1 INVX1_267 ( .A(micro_hash_synth_W_13__6_), .Y(_2504_) );
	INVX1 INVX1_268 ( .A(micro_hash_synth_W_24__6_), .Y(_2505_) );
	OAI21X1 OAI21X1_311 ( .A(_2504_), .B(micro_hash_synth_W_18__6_), .C(_2505_), .Y(_2506_) );
	AOI21X1 AOI21X1_259 ( .A(_2504_), .B(micro_hash_synth_W_18__6_), .C(_2506_), .Y(_2507_) );
	OAI22X1 OAI22X1_27 ( .A(_2503_), .B(_2471__bF_buf7), .C(_2473__bF_buf9), .D(_2507_), .Y(_1125_) );
	INVX1 INVX1_269 ( .A(micro_hash_synth_W_27__7_), .Y(_2508_) );
	INVX1 INVX1_270 ( .A(micro_hash_synth_W_13__7_), .Y(_2509_) );
	INVX1 INVX1_271 ( .A(micro_hash_synth_W_24__7_), .Y(_2510_) );
	OAI21X1 OAI21X1_312 ( .A(_2509_), .B(micro_hash_synth_W_18__7_), .C(_2510_), .Y(_2511_) );
	AOI21X1 AOI21X1_260 ( .A(_2509_), .B(micro_hash_synth_W_18__7_), .C(_2511_), .Y(_2512_) );
	OAI22X1 OAI22X1_28 ( .A(_2508_), .B(_2471__bF_buf6), .C(_2473__bF_buf8), .D(_2512_), .Y(_1136_) );
	INVX1 INVX1_272 ( .A(micro_hash_synth_W_9__0_), .Y(_2513_) );
	INVX1 INVX1_273 ( .A(bloque_in_72_), .Y(_2514_) );
	OAI22X1 OAI22X1_29 ( .A(_2513_), .B(_2471__bF_buf5), .C(_2473__bF_buf7), .D(_2514_), .Y(_1147_) );
	INVX1 INVX1_274 ( .A(micro_hash_synth_W_9__1_), .Y(_2515_) );
	INVX1 INVX1_275 ( .A(bloque_in_73_), .Y(_2516_) );
	OAI22X1 OAI22X1_30 ( .A(_2515_), .B(_2471__bF_buf4), .C(_2473__bF_buf6), .D(_2516_), .Y(_1158_) );
	INVX1 INVX1_276 ( .A(micro_hash_synth_W_9__2_), .Y(_2517_) );
	INVX1 INVX1_277 ( .A(bloque_in_74_), .Y(_2518_) );
	OAI22X1 OAI22X1_31 ( .A(_2517_), .B(_2471__bF_buf3), .C(_2473__bF_buf5), .D(_2518_), .Y(_1169_) );
	INVX1 INVX1_278 ( .A(micro_hash_synth_W_9__3_), .Y(_2519_) );
	INVX1 INVX1_279 ( .A(bloque_in_75_), .Y(_2520_) );
	OAI22X1 OAI22X1_32 ( .A(_2519_), .B(_2471__bF_buf2), .C(_2473__bF_buf4), .D(_2520_), .Y(_1176_) );
	INVX1 INVX1_280 ( .A(micro_hash_synth_W_9__4_), .Y(_2521_) );
	INVX1 INVX1_281 ( .A(bloque_in_76_), .Y(_2522_) );
	OAI22X1 OAI22X1_33 ( .A(_2521_), .B(_2471__bF_buf1), .C(_2473__bF_buf3), .D(_2522_), .Y(_1177_) );
	INVX1 INVX1_282 ( .A(micro_hash_synth_W_9__5_), .Y(_2523_) );
	INVX1 INVX1_283 ( .A(bloque_in_77_), .Y(_2524_) );
	OAI22X1 OAI22X1_34 ( .A(_2523_), .B(_2471__bF_buf0), .C(_2473__bF_buf2), .D(_2524_), .Y(_1178_) );
	INVX1 INVX1_284 ( .A(micro_hash_synth_W_9__6_), .Y(_2525_) );
	INVX1 INVX1_285 ( .A(bloque_in_78_), .Y(_2526_) );
	OAI22X1 OAI22X1_35 ( .A(_2525_), .B(_2471__bF_buf13), .C(_2473__bF_buf1), .D(_2526_), .Y(_1179_) );
	INVX1 INVX1_286 ( .A(micro_hash_synth_W_9__7_), .Y(_2527_) );
	INVX1 INVX1_287 ( .A(bloque_in_79_), .Y(_2528_) );
	OAI22X1 OAI22X1_36 ( .A(_2527_), .B(_2471__bF_buf12), .C(_2473__bF_buf0), .D(_2528_), .Y(_1180_) );
	INVX1 INVX1_288 ( .A(micro_hash_synth_W_26__0_), .Y(_2529_) );
	INVX1 INVX1_289 ( .A(micro_hash_synth_W_12__0_), .Y(_2530_) );
	INVX1 INVX1_290 ( .A(micro_hash_synth_W_23__0_), .Y(_2531_) );
	OAI21X1 OAI21X1_313 ( .A(_2530_), .B(micro_hash_synth_W_17__0_), .C(_2531_), .Y(_2532_) );
	AOI21X1 AOI21X1_261 ( .A(_2530_), .B(micro_hash_synth_W_17__0_), .C(_2532_), .Y(_2533_) );
	OAI22X1 OAI22X1_37 ( .A(_2529_), .B(_2471__bF_buf11), .C(_2473__bF_buf15), .D(_2533_), .Y(_1188_) );
	INVX1 INVX1_291 ( .A(micro_hash_synth_W_26__1_), .Y(_2534_) );
	INVX1 INVX1_292 ( .A(micro_hash_synth_W_12__1_), .Y(_2535_) );
	INVX1 INVX1_293 ( .A(micro_hash_synth_W_23__1_), .Y(_2536_) );
	OAI21X1 OAI21X1_314 ( .A(_2535_), .B(micro_hash_synth_W_17__1_), .C(_2536_), .Y(_2537_) );
	AOI21X1 AOI21X1_262 ( .A(_2535_), .B(micro_hash_synth_W_17__1_), .C(_2537_), .Y(_2538_) );
	OAI22X1 OAI22X1_38 ( .A(_2534_), .B(_2471__bF_buf10), .C(_2473__bF_buf14), .D(_2538_), .Y(_1190_) );
	INVX1 INVX1_294 ( .A(micro_hash_synth_W_26__2_), .Y(_2539_) );
	INVX1 INVX1_295 ( .A(micro_hash_synth_W_12__2_), .Y(_2540_) );
	INVX1 INVX1_296 ( .A(micro_hash_synth_W_23__2_), .Y(_2541_) );
	OAI21X1 OAI21X1_315 ( .A(_2540_), .B(micro_hash_synth_W_17__2_), .C(_2541_), .Y(_2542_) );
	AOI21X1 AOI21X1_263 ( .A(_2540_), .B(micro_hash_synth_W_17__2_), .C(_2542_), .Y(_2543_) );
	OAI22X1 OAI22X1_39 ( .A(_2539_), .B(_2471__bF_buf9), .C(_2473__bF_buf13), .D(_2543_), .Y(_935_) );
	INVX1 INVX1_297 ( .A(micro_hash_synth_W_26__3_), .Y(_2544_) );
	INVX1 INVX1_298 ( .A(micro_hash_synth_W_12__3_), .Y(_2545_) );
	INVX1 INVX1_299 ( .A(micro_hash_synth_W_23__3_), .Y(_2546_) );
	OAI21X1 OAI21X1_316 ( .A(_2545_), .B(micro_hash_synth_W_17__3_), .C(_2546_), .Y(_2547_) );
	AOI21X1 AOI21X1_264 ( .A(_2545_), .B(micro_hash_synth_W_17__3_), .C(_2547_), .Y(_2548_) );
	OAI22X1 OAI22X1_40 ( .A(_2544_), .B(_2471__bF_buf8), .C(_2473__bF_buf12), .D(_2548_), .Y(_936_) );
	INVX1 INVX1_300 ( .A(micro_hash_synth_W_26__4_), .Y(_2549_) );
	INVX1 INVX1_301 ( .A(micro_hash_synth_W_12__4_), .Y(_2550_) );
	INVX1 INVX1_302 ( .A(micro_hash_synth_W_23__4_), .Y(_2551_) );
	OAI21X1 OAI21X1_317 ( .A(_2550_), .B(micro_hash_synth_W_17__4_), .C(_2551_), .Y(_2552_) );
	AOI21X1 AOI21X1_265 ( .A(_2550_), .B(micro_hash_synth_W_17__4_), .C(_2552_), .Y(_2553_) );
	OAI22X1 OAI22X1_41 ( .A(_2549_), .B(_2471__bF_buf7), .C(_2473__bF_buf11), .D(_2553_), .Y(_937_) );
	INVX1 INVX1_303 ( .A(micro_hash_synth_W_26__5_), .Y(_2554_) );
	INVX1 INVX1_304 ( .A(micro_hash_synth_W_12__5_), .Y(_2555_) );
	INVX1 INVX1_305 ( .A(micro_hash_synth_W_23__5_), .Y(_2556_) );
	OAI21X1 OAI21X1_318 ( .A(_2555_), .B(micro_hash_synth_W_17__5_), .C(_2556_), .Y(_2557_) );
	AOI21X1 AOI21X1_266 ( .A(_2555_), .B(micro_hash_synth_W_17__5_), .C(_2557_), .Y(_2558_) );
	OAI22X1 OAI22X1_42 ( .A(_2554_), .B(_2471__bF_buf6), .C(_2473__bF_buf10), .D(_2558_), .Y(_938_) );
	INVX1 INVX1_306 ( .A(micro_hash_synth_W_26__6_), .Y(_2559_) );
	INVX1 INVX1_307 ( .A(micro_hash_synth_W_12__6_), .Y(_2560_) );
	INVX1 INVX1_308 ( .A(micro_hash_synth_W_23__6_), .Y(_2561_) );
	OAI21X1 OAI21X1_319 ( .A(_2560_), .B(micro_hash_synth_W_17__6_), .C(_2561_), .Y(_2562_) );
	AOI21X1 AOI21X1_267 ( .A(_2560_), .B(micro_hash_synth_W_17__6_), .C(_2562_), .Y(_2563_) );
	OAI22X1 OAI22X1_43 ( .A(_2559_), .B(_2471__bF_buf5), .C(_2473__bF_buf9), .D(_2563_), .Y(_939_) );
	INVX1 INVX1_309 ( .A(micro_hash_synth_W_26__7_), .Y(_2564_) );
	INVX1 INVX1_310 ( .A(micro_hash_synth_W_12__7_), .Y(_2565_) );
	INVX1 INVX1_311 ( .A(micro_hash_synth_W_23__7_), .Y(_2566_) );
	OAI21X1 OAI21X1_320 ( .A(_2565_), .B(micro_hash_synth_W_17__7_), .C(_2566_), .Y(_2567_) );
	AOI21X1 AOI21X1_268 ( .A(_2565_), .B(micro_hash_synth_W_17__7_), .C(_2567_), .Y(_2568_) );
	OAI22X1 OAI22X1_44 ( .A(_2564_), .B(_2471__bF_buf4), .C(_2473__bF_buf8), .D(_2568_), .Y(_940_) );
	INVX1 INVX1_312 ( .A(micro_hash_synth_W_25__0_), .Y(_2569_) );
	INVX1 INVX1_313 ( .A(micro_hash_synth_W_11__0_), .Y(_2570_) );
	INVX1 INVX1_314 ( .A(micro_hash_synth_W_22__0_), .Y(_2571_) );
	OAI21X1 OAI21X1_321 ( .A(_2570_), .B(micro_hash_synth_W_16__0_), .C(_2571_), .Y(_2572_) );
	AOI21X1 AOI21X1_269 ( .A(_2570_), .B(micro_hash_synth_W_16__0_), .C(_2572_), .Y(_2573_) );
	OAI22X1 OAI22X1_45 ( .A(_2569_), .B(_2471__bF_buf3), .C(_2473__bF_buf7), .D(_2573_), .Y(_941_) );
	INVX1 INVX1_315 ( .A(micro_hash_synth_W_25__1_), .Y(_2574_) );
	INVX1 INVX1_316 ( .A(micro_hash_synth_W_11__1_), .Y(_2575_) );
	INVX1 INVX1_317 ( .A(micro_hash_synth_W_22__1_), .Y(_2576_) );
	OAI21X1 OAI21X1_322 ( .A(_2575_), .B(micro_hash_synth_W_16__1_), .C(_2576_), .Y(_2577_) );
	AOI21X1 AOI21X1_270 ( .A(_2575_), .B(micro_hash_synth_W_16__1_), .C(_2577_), .Y(_2578_) );
	OAI22X1 OAI22X1_46 ( .A(_2574_), .B(_2471__bF_buf2), .C(_2473__bF_buf6), .D(_2578_), .Y(_950_) );
	INVX1 INVX1_318 ( .A(micro_hash_synth_W_25__2_), .Y(_2579_) );
	INVX1 INVX1_319 ( .A(micro_hash_synth_W_11__2_), .Y(_2580_) );
	INVX1 INVX1_320 ( .A(micro_hash_synth_W_22__2_), .Y(_2581_) );
	OAI21X1 OAI21X1_323 ( .A(_2580_), .B(micro_hash_synth_W_16__2_), .C(_2581_), .Y(_2582_) );
	AOI21X1 AOI21X1_271 ( .A(_2580_), .B(micro_hash_synth_W_16__2_), .C(_2582_), .Y(_2583_) );
	OAI22X1 OAI22X1_47 ( .A(_2579_), .B(_2471__bF_buf1), .C(_2473__bF_buf5), .D(_2583_), .Y(_955_) );
	INVX1 INVX1_321 ( .A(micro_hash_synth_W_25__3_), .Y(_2584_) );
	INVX1 INVX1_322 ( .A(micro_hash_synth_W_11__3_), .Y(_2585_) );
	INVX1 INVX1_323 ( .A(micro_hash_synth_W_22__3_), .Y(_2586_) );
	OAI21X1 OAI21X1_324 ( .A(_2585_), .B(micro_hash_synth_W_16__3_), .C(_2586_), .Y(_2587_) );
	AOI21X1 AOI21X1_272 ( .A(_2585_), .B(micro_hash_synth_W_16__3_), .C(_2587_), .Y(_2588_) );
	OAI22X1 OAI22X1_48 ( .A(_2584_), .B(_2471__bF_buf0), .C(_2473__bF_buf4), .D(_2588_), .Y(_971_) );
	INVX1 INVX1_324 ( .A(micro_hash_synth_W_25__4_), .Y(_2589_) );
	INVX1 INVX1_325 ( .A(micro_hash_synth_W_11__4_), .Y(_2590_) );
	INVX1 INVX1_326 ( .A(micro_hash_synth_W_22__4_), .Y(_2591_) );
	OAI21X1 OAI21X1_325 ( .A(_2590_), .B(micro_hash_synth_W_16__4_), .C(_2591_), .Y(_2592_) );
	AOI21X1 AOI21X1_273 ( .A(_2590_), .B(micro_hash_synth_W_16__4_), .C(_2592_), .Y(_2593_) );
	OAI22X1 OAI22X1_49 ( .A(_2589_), .B(_2471__bF_buf13), .C(_2473__bF_buf3), .D(_2593_), .Y(_987_) );
	INVX1 INVX1_327 ( .A(micro_hash_synth_W_25__5_), .Y(_2594_) );
	INVX1 INVX1_328 ( .A(micro_hash_synth_W_11__5_), .Y(_2595_) );
	INVX1 INVX1_329 ( .A(micro_hash_synth_W_22__5_), .Y(_2596_) );
	OAI21X1 OAI21X1_326 ( .A(_2595_), .B(micro_hash_synth_W_16__5_), .C(_2596_), .Y(_2597_) );
	AOI21X1 AOI21X1_274 ( .A(_2595_), .B(micro_hash_synth_W_16__5_), .C(_2597_), .Y(_2598_) );
	OAI22X1 OAI22X1_50 ( .A(_2594_), .B(_2471__bF_buf12), .C(_2473__bF_buf2), .D(_2598_), .Y(_1003_) );
	INVX1 INVX1_330 ( .A(micro_hash_synth_W_25__6_), .Y(_2599_) );
	INVX1 INVX1_331 ( .A(micro_hash_synth_W_11__6_), .Y(_2600_) );
	INVX1 INVX1_332 ( .A(micro_hash_synth_W_22__6_), .Y(_2601_) );
	OAI21X1 OAI21X1_327 ( .A(_2600_), .B(micro_hash_synth_W_16__6_), .C(_2601_), .Y(_2602_) );
	AOI21X1 AOI21X1_275 ( .A(_2600_), .B(micro_hash_synth_W_16__6_), .C(_2602_), .Y(_2603_) );
	OAI22X1 OAI22X1_51 ( .A(_2599_), .B(_2471__bF_buf11), .C(_2473__bF_buf1), .D(_2603_), .Y(_1019_) );
	INVX1 INVX1_333 ( .A(micro_hash_synth_W_25__7_), .Y(_2604_) );
	INVX1 INVX1_334 ( .A(micro_hash_synth_W_11__7_), .Y(_2605_) );
	INVX1 INVX1_335 ( .A(micro_hash_synth_W_22__7_), .Y(_2606_) );
	OAI21X1 OAI21X1_328 ( .A(_2605_), .B(micro_hash_synth_W_16__7_), .C(_2606_), .Y(_2607_) );
	AOI21X1 AOI21X1_276 ( .A(_2605_), .B(micro_hash_synth_W_16__7_), .C(_2607_), .Y(_2608_) );
	OAI22X1 OAI22X1_52 ( .A(_2604_), .B(_2471__bF_buf10), .C(_2473__bF_buf0), .D(_2608_), .Y(_1035_) );
	NOR2X1 NOR2X1_94 ( .A(concatenador_count_0_bF_buf8), .B(_2463_), .Y(_2609_) );
	INVX1 INVX1_336 ( .A(concatenador_count_5_), .Y(_2610_) );
	NOR2X1 NOR2X1_95 ( .A(_1__bF_buf5), .B(_2610_), .Y(_2611_) );
	AND2X2 AND2X2_23 ( .A(_2609__bF_buf3), .B(_2611_), .Y(_2612_) );
	NAND2X1 NAND2X1_106 ( .A(_2466_), .B(_2612_), .Y(_2613_) );
	OAI21X1 OAI21X1_329 ( .A(_2467_), .B(concatenador_count_5_), .C(H_16_), .Y(_1191_) );
	AND2X2 AND2X2_24 ( .A(H_16_), .B(micro_hash_synth_c_0_), .Y(_1192_) );
	NOR2X1 NOR2X1_96 ( .A(H_16_), .B(micro_hash_synth_c_0_), .Y(_1193_) );
	NOR2X1 NOR2X1_97 ( .A(_1193_), .B(_1192_), .Y(_1194_) );
	OAI21X1 OAI21X1_330 ( .A(_2613_), .B(_1194_), .C(reset_L_bF_buf3), .Y(_1195_) );
	AOI21X1 AOI21X1_277 ( .A(_2613_), .B(_1191_), .C(_1195_), .Y(_927__16_) );
	INVX4 INVX4_4 ( .A(_2613_), .Y(_1196_) );
	XOR2X1 XOR2X1_12 ( .A(H_17_), .B(micro_hash_synth_c_1_), .Y(_1197_) );
	NAND2X1 NAND2X1_107 ( .A(_1192_), .B(_1197_), .Y(_1198_) );
	OR2X2 OR2X2_22 ( .A(_1197_), .B(_1192_), .Y(_1199_) );
	NAND3X1 NAND3X1_74 ( .A(_1198_), .B(_1199_), .C(_1196__bF_buf3), .Y(_1200_) );
	OAI21X1 OAI21X1_331 ( .A(_2468_), .B(H_17_), .C(_2613_), .Y(_1201_) );
	NAND3X1 NAND3X1_75 ( .A(reset_L_bF_buf2), .B(_1200_), .C(_1201_), .Y(_927__17_) );
	INVX8 INVX8_3 ( .A(reset_L_bF_buf1), .Y(_1202_) );
	NOR2X1 NOR2X1_98 ( .A(_1202__bF_buf5), .B(_2613_), .Y(_1203_) );
	INVX4 INVX4_5 ( .A(_1203_), .Y(_1204_) );
	OAI21X1 OAI21X1_332 ( .A(_2467_), .B(concatenador_count_5_), .C(reset_L_bF_buf0), .Y(_1205_) );
	OAI21X1 OAI21X1_333 ( .A(_1205__bF_buf3), .B(H_18_), .C(_1204_), .Y(_1206_) );
	INVX1 INVX1_337 ( .A(H_17_), .Y(_1207_) );
	INVX1 INVX1_338 ( .A(micro_hash_synth_c_1_), .Y(_1208_) );
	OAI21X1 OAI21X1_334 ( .A(_1207_), .B(_1208_), .C(_1198_), .Y(_1209_) );
	XOR2X1 XOR2X1_13 ( .A(H_18_), .B(micro_hash_synth_c_2_), .Y(_1210_) );
	NAND2X1 NAND2X1_108 ( .A(_1210_), .B(_1209_), .Y(_1211_) );
	INVX1 INVX1_339 ( .A(_1211_), .Y(_1212_) );
	OAI21X1 OAI21X1_335 ( .A(_1209_), .B(_1210_), .C(_1196__bF_buf2), .Y(_1213_) );
	OAI21X1 OAI21X1_336 ( .A(_1212_), .B(_1213_), .C(_1206_), .Y(_927__18_) );
	OAI21X1 OAI21X1_337 ( .A(_1205__bF_buf2), .B(H_19_), .C(_1204_), .Y(_1214_) );
	INVX1 INVX1_340 ( .A(H_18_), .Y(_1215_) );
	INVX1 INVX1_341 ( .A(micro_hash_synth_c_2_), .Y(_1216_) );
	OAI21X1 OAI21X1_338 ( .A(_1215_), .B(_1216_), .C(_1211_), .Y(_1217_) );
	NOR2X1 NOR2X1_99 ( .A(H_19_), .B(micro_hash_synth_c_3_), .Y(_1218_) );
	NAND2X1 NAND2X1_109 ( .A(H_19_), .B(micro_hash_synth_c_3_), .Y(_1219_) );
	INVX1 INVX1_342 ( .A(_1219_), .Y(_1220_) );
	NOR2X1 NOR2X1_100 ( .A(_1218_), .B(_1220_), .Y(_1221_) );
	AND2X2 AND2X2_25 ( .A(_1217_), .B(_1221_), .Y(_1222_) );
	OAI21X1 OAI21X1_339 ( .A(_1217_), .B(_1221_), .C(_1196__bF_buf1), .Y(_1223_) );
	OAI21X1 OAI21X1_340 ( .A(_1222_), .B(_1223_), .C(_1214_), .Y(_927__19_) );
	OAI21X1 OAI21X1_341 ( .A(_1205__bF_buf1), .B(H_20_), .C(_1204_), .Y(_1224_) );
	XOR2X1 XOR2X1_14 ( .A(H_20_), .B(micro_hash_synth_c_4_), .Y(_1225_) );
	INVX1 INVX1_343 ( .A(_1225_), .Y(_1226_) );
	INVX1 INVX1_344 ( .A(_1218_), .Y(_1227_) );
	AOI21X1 AOI21X1_278 ( .A(_1227_), .B(_1217_), .C(_1220_), .Y(_1228_) );
	NAND2X1 NAND2X1_110 ( .A(_1226_), .B(_1228_), .Y(_1229_) );
	INVX1 INVX1_345 ( .A(_1229_), .Y(_1230_) );
	OAI21X1 OAI21X1_342 ( .A(_1228_), .B(_1226_), .C(_1196__bF_buf0), .Y(_1231_) );
	OAI21X1 OAI21X1_343 ( .A(_1230_), .B(_1231_), .C(_1224_), .Y(_927__20_) );
	OAI21X1 OAI21X1_344 ( .A(_1205__bF_buf0), .B(H_21_), .C(_1204_), .Y(_1232_) );
	NAND2X1 NAND2X1_111 ( .A(H_20_), .B(micro_hash_synth_c_4_), .Y(_1233_) );
	OAI21X1 OAI21X1_345 ( .A(_1228_), .B(_1226_), .C(_1233_), .Y(_1234_) );
	XOR2X1 XOR2X1_15 ( .A(H_21_), .B(micro_hash_synth_c_5_), .Y(_1235_) );
	AND2X2 AND2X2_26 ( .A(_1234_), .B(_1235_), .Y(_1236_) );
	OAI21X1 OAI21X1_346 ( .A(_1234_), .B(_1235_), .C(_1196__bF_buf3), .Y(_1237_) );
	OAI21X1 OAI21X1_347 ( .A(_1236_), .B(_1237_), .C(_1232_), .Y(_927__21_) );
	OAI21X1 OAI21X1_348 ( .A(_1205__bF_buf3), .B(H_22_), .C(_1204_), .Y(_1238_) );
	XOR2X1 XOR2X1_16 ( .A(H_22_), .B(micro_hash_synth_c_6_), .Y(_1239_) );
	NAND2X1 NAND2X1_112 ( .A(H_21_), .B(micro_hash_synth_c_5_), .Y(_1240_) );
	OAI21X1 OAI21X1_349 ( .A(H_21_), .B(micro_hash_synth_c_5_), .C(_1234_), .Y(_1241_) );
	NAND2X1 NAND2X1_113 ( .A(_1240_), .B(_1241_), .Y(_1242_) );
	NOR2X1 NOR2X1_101 ( .A(_1239_), .B(_1242_), .Y(_1243_) );
	NAND2X1 NAND2X1_114 ( .A(_1239_), .B(_1242_), .Y(_1244_) );
	NAND2X1 NAND2X1_115 ( .A(_1196__bF_buf2), .B(_1244_), .Y(_1245_) );
	OAI21X1 OAI21X1_350 ( .A(_1245_), .B(_1243_), .C(_1238_), .Y(_927__22_) );
	NAND2X1 NAND2X1_116 ( .A(H_22_), .B(micro_hash_synth_c_6_), .Y(_1246_) );
	NAND2X1 NAND2X1_117 ( .A(_1246_), .B(_1244_), .Y(_1247_) );
	XOR2X1 XOR2X1_17 ( .A(H_23_), .B(micro_hash_synth_c_7_), .Y(_1248_) );
	AND2X2 AND2X2_27 ( .A(_1247_), .B(_1248_), .Y(_1249_) );
	OAI21X1 OAI21X1_351 ( .A(_1247_), .B(_1248_), .C(_1196__bF_buf1), .Y(_1250_) );
	OAI21X1 OAI21X1_352 ( .A(_1205__bF_buf2), .B(H_23_), .C(_1204_), .Y(_1251_) );
	OAI21X1 OAI21X1_353 ( .A(_1249_), .B(_1250_), .C(_1251_), .Y(_927__23_) );
	INVX1 INVX1_346 ( .A(H_8_), .Y(_1252_) );
	NOR2X1 NOR2X1_102 ( .A(_1202__bF_buf4), .B(_1196__bF_buf0), .Y(_1253_) );
	INVX2 INVX2_2 ( .A(_1253_), .Y(_1254_) );
	OAI22X1 OAI22X1_53 ( .A(micro_hash_synth_b_0_), .B(_1204_), .C(_1254_), .D(_2468_), .Y(_1255_) );
	INVX1 INVX1_347 ( .A(micro_hash_synth_b_0_), .Y(_1256_) );
	NOR2X1 NOR2X1_103 ( .A(_1252_), .B(_1256_), .Y(_1257_) );
	AOI22X1 AOI22X1_24 ( .A(_1203_), .B(_1257_), .C(_1255_), .D(_1252_), .Y(_927__8_) );
	XOR2X1 XOR2X1_18 ( .A(H_9_), .B(micro_hash_synth_b_1_), .Y(_1258_) );
	XNOR2X1 XNOR2X1_13 ( .A(_1258_), .B(_1257_), .Y(_1259_) );
	OAI21X1 OAI21X1_354 ( .A(_2467_), .B(concatenador_count_5_), .C(H_9_), .Y(_1260_) );
	OAI22X1 OAI22X1_54 ( .A(_1204_), .B(_1259_), .C(_1254_), .D(_1260_), .Y(_927__9_) );
	INVX1 INVX1_348 ( .A(H_9_), .Y(_1261_) );
	INVX1 INVX1_349 ( .A(micro_hash_synth_b_1_), .Y(_1262_) );
	NAND2X1 NAND2X1_118 ( .A(_1257_), .B(_1258_), .Y(_1263_) );
	OAI21X1 OAI21X1_355 ( .A(_1261_), .B(_1262_), .C(_1263_), .Y(_1264_) );
	NOR2X1 NOR2X1_104 ( .A(H_10_), .B(micro_hash_synth_b_2_), .Y(_1265_) );
	AND2X2 AND2X2_28 ( .A(H_10_), .B(micro_hash_synth_b_2_), .Y(_1266_) );
	NOR2X1 NOR2X1_105 ( .A(_1265_), .B(_1266_), .Y(_1267_) );
	XNOR2X1 XNOR2X1_14 ( .A(_1264_), .B(_1267_), .Y(_1268_) );
	INVX4 INVX4_6 ( .A(_1205__bF_buf1), .Y(_1269_) );
	NAND2X1 NAND2X1_119 ( .A(H_10_), .B(_1269__bF_buf3), .Y(_1270_) );
	AOI22X1 AOI22X1_25 ( .A(_1196__bF_buf3), .B(_1268_), .C(_1270_), .D(_1204_), .Y(_927__10_) );
	OAI21X1 OAI21X1_356 ( .A(_1205__bF_buf0), .B(H_11_), .C(_1204_), .Y(_1271_) );
	AOI21X1 AOI21X1_279 ( .A(_1267_), .B(_1264_), .C(_1266_), .Y(_1272_) );
	NOR2X1 NOR2X1_106 ( .A(H_11_), .B(micro_hash_synth_b_3_), .Y(_1273_) );
	NAND2X1 NAND2X1_120 ( .A(H_11_), .B(micro_hash_synth_b_3_), .Y(_1274_) );
	INVX1 INVX1_350 ( .A(_1274_), .Y(_1275_) );
	NOR2X1 NOR2X1_107 ( .A(_1273_), .B(_1275_), .Y(_1276_) );
	INVX1 INVX1_351 ( .A(_1276_), .Y(_1277_) );
	AND2X2 AND2X2_29 ( .A(_1272_), .B(_1277_), .Y(_1278_) );
	OAI21X1 OAI21X1_357 ( .A(_1272_), .B(_1277_), .C(_1196__bF_buf2), .Y(_1279_) );
	OAI21X1 OAI21X1_358 ( .A(_1278_), .B(_1279_), .C(_1271_), .Y(_927__11_) );
	XOR2X1 XOR2X1_19 ( .A(H_12_), .B(micro_hash_synth_b_4_), .Y(_1280_) );
	OAI21X1 OAI21X1_359 ( .A(_1272_), .B(_1273_), .C(_1274_), .Y(_1281_) );
	XNOR2X1 XNOR2X1_15 ( .A(_1281_), .B(_1280_), .Y(_1282_) );
	AOI21X1 AOI21X1_280 ( .A(H_12_), .B(_1269__bF_buf2), .C(_1203_), .Y(_1283_) );
	AOI21X1 AOI21X1_281 ( .A(_1196__bF_buf1), .B(_1282_), .C(_1283_), .Y(_927__12_) );
	AOI21X1 AOI21X1_282 ( .A(H_13_), .B(_1269__bF_buf1), .C(_1203_), .Y(_1284_) );
	AND2X2 AND2X2_30 ( .A(H_12_), .B(micro_hash_synth_b_4_), .Y(_1285_) );
	AOI21X1 AOI21X1_283 ( .A(_1280_), .B(_1281_), .C(_1285_), .Y(_1286_) );
	NOR2X1 NOR2X1_108 ( .A(H_13_), .B(micro_hash_synth_b_5_), .Y(_1287_) );
	NAND2X1 NAND2X1_121 ( .A(H_13_), .B(micro_hash_synth_b_5_), .Y(_1288_) );
	INVX1 INVX1_352 ( .A(_1288_), .Y(_1289_) );
	NOR2X1 NOR2X1_109 ( .A(_1287_), .B(_1289_), .Y(_1290_) );
	XOR2X1 XOR2X1_20 ( .A(_1286_), .B(_1290_), .Y(_1291_) );
	AOI21X1 AOI21X1_284 ( .A(_1196__bF_buf0), .B(_1291_), .C(_1284_), .Y(_927__13_) );
	XOR2X1 XOR2X1_21 ( .A(H_14_), .B(micro_hash_synth_b_6_), .Y(_1292_) );
	OAI21X1 OAI21X1_360 ( .A(_1286_), .B(_1287_), .C(_1288_), .Y(_1293_) );
	XNOR2X1 XNOR2X1_16 ( .A(_1293_), .B(_1292_), .Y(_1294_) );
	AOI21X1 AOI21X1_285 ( .A(H_14_), .B(_1269__bF_buf0), .C(_1203_), .Y(_1295_) );
	AOI21X1 AOI21X1_286 ( .A(_1196__bF_buf3), .B(_1294_), .C(_1295_), .Y(_927__14_) );
	NAND2X1 NAND2X1_122 ( .A(H_14_), .B(micro_hash_synth_b_6_), .Y(_1296_) );
	NAND2X1 NAND2X1_123 ( .A(_1292_), .B(_1293_), .Y(_1297_) );
	XNOR2X1 XNOR2X1_17 ( .A(H_15_), .B(micro_hash_synth_b_7_), .Y(_1298_) );
	AOI21X1 AOI21X1_287 ( .A(_1296_), .B(_1297_), .C(_1298_), .Y(_1299_) );
	NAND2X1 NAND2X1_124 ( .A(_1296_), .B(_1297_), .Y(_1300_) );
	INVX1 INVX1_353 ( .A(_1298_), .Y(_1301_) );
	OAI21X1 OAI21X1_361 ( .A(_1300_), .B(_1301_), .C(_1196__bF_buf2), .Y(_1302_) );
	OAI21X1 OAI21X1_362 ( .A(_1205__bF_buf3), .B(H_15_), .C(_1204_), .Y(_1303_) );
	OAI21X1 OAI21X1_363 ( .A(_1302_), .B(_1299_), .C(_1303_), .Y(_927__15_) );
	INVX1 INVX1_354 ( .A(H_0_), .Y(_1304_) );
	OAI22X1 OAI22X1_55 ( .A(micro_hash_synth_a_0_), .B(_1204_), .C(_1254_), .D(_2468_), .Y(_1305_) );
	INVX1 INVX1_355 ( .A(micro_hash_synth_a_0_), .Y(_1306_) );
	NOR2X1 NOR2X1_110 ( .A(_1304_), .B(_1306_), .Y(_1307_) );
	AOI22X1 AOI22X1_26 ( .A(_1203_), .B(_1307_), .C(_1305_), .D(_1304_), .Y(_927__0_) );
	NOR2X1 NOR2X1_111 ( .A(H_1_), .B(micro_hash_synth_a_1_), .Y(_1308_) );
	INVX1 INVX1_356 ( .A(H_1_), .Y(_1309_) );
	INVX1 INVX1_357 ( .A(micro_hash_synth_a_1_), .Y(_1310_) );
	NOR2X1 NOR2X1_112 ( .A(_1309_), .B(_1310_), .Y(_1311_) );
	NOR2X1 NOR2X1_113 ( .A(_1308_), .B(_1311_), .Y(_1312_) );
	NAND2X1 NAND2X1_125 ( .A(_1307_), .B(_1312_), .Y(_1313_) );
	OR2X2 OR2X2_23 ( .A(_1312_), .B(_1307_), .Y(_1314_) );
	AOI21X1 AOI21X1_288 ( .A(_1313_), .B(_1314_), .C(_2613_), .Y(_1315_) );
	NAND2X1 NAND2X1_126 ( .A(H_1_), .B(_1269__bF_buf3), .Y(_1316_) );
	AOI21X1 AOI21X1_289 ( .A(_1204_), .B(_1316_), .C(_1315_), .Y(_927__1_) );
	OAI21X1 OAI21X1_364 ( .A(_1309_), .B(_1310_), .C(_1313_), .Y(_1317_) );
	NOR2X1 NOR2X1_114 ( .A(H_2_), .B(micro_hash_synth_a_2_), .Y(_1318_) );
	AND2X2 AND2X2_31 ( .A(H_2_), .B(micro_hash_synth_a_2_), .Y(_1319_) );
	NOR2X1 NOR2X1_115 ( .A(_1318_), .B(_1319_), .Y(_1320_) );
	XNOR2X1 XNOR2X1_18 ( .A(_1317_), .B(_1320_), .Y(_1321_) );
	NAND2X1 NAND2X1_127 ( .A(H_2_), .B(_1269__bF_buf2), .Y(_1322_) );
	AOI22X1 AOI22X1_27 ( .A(_1196__bF_buf1), .B(_1321_), .C(_1322_), .D(_1204_), .Y(_927__2_) );
	AOI21X1 AOI21X1_290 ( .A(H_3_), .B(_1269__bF_buf1), .C(_1203_), .Y(_1323_) );
	AOI21X1 AOI21X1_291 ( .A(_1320_), .B(_1317_), .C(_1319_), .Y(_1324_) );
	NOR2X1 NOR2X1_116 ( .A(H_3_), .B(micro_hash_synth_a_3_), .Y(_1325_) );
	INVX1 INVX1_358 ( .A(_1325_), .Y(_1326_) );
	NAND2X1 NAND2X1_128 ( .A(H_3_), .B(micro_hash_synth_a_3_), .Y(_1327_) );
	NAND2X1 NAND2X1_129 ( .A(_1327_), .B(_1326_), .Y(_1328_) );
	XNOR2X1 XNOR2X1_19 ( .A(_1324_), .B(_1328_), .Y(_1329_) );
	AOI21X1 AOI21X1_292 ( .A(_1196__bF_buf0), .B(_1329_), .C(_1323_), .Y(_927__3_) );
	XOR2X1 XOR2X1_22 ( .A(H_4_), .B(micro_hash_synth_a_4_), .Y(_1330_) );
	OAI21X1 OAI21X1_365 ( .A(_1324_), .B(_1325_), .C(_1327_), .Y(_1331_) );
	XNOR2X1 XNOR2X1_20 ( .A(_1331_), .B(_1330_), .Y(_1332_) );
	AOI21X1 AOI21X1_293 ( .A(H_4_), .B(_1269__bF_buf0), .C(_1203_), .Y(_1333_) );
	AOI21X1 AOI21X1_294 ( .A(_1196__bF_buf3), .B(_1332_), .C(_1333_), .Y(_927__4_) );
	AOI21X1 AOI21X1_295 ( .A(H_5_), .B(_1269__bF_buf3), .C(_1203_), .Y(_1334_) );
	AND2X2 AND2X2_32 ( .A(H_4_), .B(micro_hash_synth_a_4_), .Y(_1335_) );
	AOI21X1 AOI21X1_296 ( .A(_1330_), .B(_1331_), .C(_1335_), .Y(_1336_) );
	NOR2X1 NOR2X1_117 ( .A(H_5_), .B(micro_hash_synth_a_5_), .Y(_1337_) );
	NAND2X1 NAND2X1_130 ( .A(H_5_), .B(micro_hash_synth_a_5_), .Y(_1338_) );
	INVX1 INVX1_359 ( .A(_1338_), .Y(_1339_) );
	NOR2X1 NOR2X1_118 ( .A(_1337_), .B(_1339_), .Y(_1340_) );
	OAI21X1 OAI21X1_366 ( .A(_1336_), .B(_1340_), .C(_1196__bF_buf2), .Y(_1341_) );
	AOI21X1 AOI21X1_297 ( .A(_1336_), .B(_1340_), .C(_1341_), .Y(_1342_) );
	NOR2X1 NOR2X1_119 ( .A(_1334_), .B(_1342_), .Y(_927__5_) );
	XOR2X1 XOR2X1_23 ( .A(H_6_), .B(micro_hash_synth_a_6_), .Y(_1343_) );
	OAI21X1 OAI21X1_367 ( .A(_1336_), .B(_1337_), .C(_1338_), .Y(_1344_) );
	XNOR2X1 XNOR2X1_21 ( .A(_1344_), .B(_1343_), .Y(_1345_) );
	AOI21X1 AOI21X1_298 ( .A(H_6_), .B(_1269__bF_buf2), .C(_1203_), .Y(_1346_) );
	AOI21X1 AOI21X1_299 ( .A(_1196__bF_buf1), .B(_1345_), .C(_1346_), .Y(_927__6_) );
	AOI21X1 AOI21X1_300 ( .A(H_7_), .B(_1269__bF_buf1), .C(_1203_), .Y(_1347_) );
	INVX1 INVX1_360 ( .A(H_6_), .Y(_1348_) );
	INVX1 INVX1_361 ( .A(micro_hash_synth_a_6_), .Y(_1349_) );
	NAND2X1 NAND2X1_131 ( .A(_1343_), .B(_1344_), .Y(_1350_) );
	OAI21X1 OAI21X1_368 ( .A(_1348_), .B(_1349_), .C(_1350_), .Y(_1351_) );
	XOR2X1 XOR2X1_24 ( .A(H_7_), .B(micro_hash_synth_a_7_), .Y(_1352_) );
	XNOR2X1 XNOR2X1_22 ( .A(_1351_), .B(_1352_), .Y(_1353_) );
	AOI21X1 AOI21X1_301 ( .A(_1196__bF_buf0), .B(_1353_), .C(_1347_), .Y(_927__7_) );
	NAND2X1 NAND2X1_132 ( .A(concatenador_count_5_), .B(_2467_), .Y(_1354_) );
	NOR2X1 NOR2X1_120 ( .A(_1202__bF_buf3), .B(_1354__bF_buf3), .Y(_1355_) );
	INVX2 INVX2_3 ( .A(_1355_), .Y(_1356_) );
	OR2X2 OR2X2_24 ( .A(_1356_), .B(micro_hash_synth_k_0_), .Y(_932__0_) );
	INVX1 INVX1_362 ( .A(micro_hash_synth_k_1_), .Y(_1357_) );
	NOR2X1 NOR2X1_121 ( .A(_1357_), .B(_1356_), .Y(_932__1_) );
	INVX1 INVX1_363 ( .A(micro_hash_synth_k_2_), .Y(_1358_) );
	NOR2X1 NOR2X1_122 ( .A(_1358_), .B(_1356_), .Y(_932__2_) );
	INVX1 INVX1_364 ( .A(micro_hash_synth_k_3_), .Y(_1359_) );
	INVX1 INVX1_365 ( .A(concatenador_count_4_), .Y(_1360_) );
	AOI21X1 AOI21X1_302 ( .A(_2464_), .B(_2470__bF_buf1), .C(_1360_), .Y(_1361_) );
	OAI21X1 OAI21X1_369 ( .A(_1361_), .B(concatenador_count_5_), .C(reset_L_bF_buf11), .Y(_1362_) );
	INVX1 INVX1_366 ( .A(_1362_), .Y(_1363_) );
	OAI21X1 OAI21X1_370 ( .A(_1354__bF_buf2), .B(_1359_), .C(_1363_), .Y(_932__3_) );
	INVX1 INVX1_367 ( .A(micro_hash_synth_k_4_), .Y(_1364_) );
	OAI21X1 OAI21X1_371 ( .A(_1354__bF_buf1), .B(_1364_), .C(_1363_), .Y(_932__4_) );
	INVX1 INVX1_368 ( .A(micro_hash_synth_k_5_), .Y(_1365_) );
	INVX4 INVX4_7 ( .A(_1354__bF_buf0), .Y(_1366_) );
	AOI21X1 AOI21X1_303 ( .A(_1365_), .B(_1366_), .C(_1362_), .Y(_932__5_) );
	AND2X2 AND2X2_33 ( .A(_1355_), .B(micro_hash_synth_k_6_), .Y(_932__6_) );
	OR2X2 OR2X2_25 ( .A(_1356_), .B(micro_hash_synth_k_7_), .Y(_932__7_) );
	INVX1 INVX1_369 ( .A(micro_hash_synth_c_0_), .Y(_1367_) );
	XOR2X1 XOR2X1_25 ( .A(micro_hash_synth_k_0_), .B(micro_hash_synth_x_0_), .Y(_1368_) );
	INVX1 INVX1_370 ( .A(_1368_), .Y(_1369_) );
	NAND2X1 NAND2X1_133 ( .A(_2463_), .B(_2464_), .Y(_1370_) );
	XNOR2X1 XNOR2X1_23 ( .A(_1370_), .B(concatenador_count_4_), .Y(_1371_) );
	INVX4 INVX4_8 ( .A(_1371_), .Y(_1372_) );
	XOR2X1 XOR2X1_26 ( .A(concatenador_count_1_bF_buf3), .B(concatenador_count_2_), .Y(_1373_) );
	MUX2X1 MUX2X1_1 ( .A(micro_hash_synth_W_29__0_), .B(micro_hash_synth_W_28__0_), .S(concatenador_count_0_bF_buf7), .Y(_1374_) );
	MUX2X1 MUX2X1_2 ( .A(micro_hash_synth_W_31__0_), .B(micro_hash_synth_W_30__0_), .S(concatenador_count_0_bF_buf6), .Y(_1375_) );
	MUX2X1 MUX2X1_3 ( .A(_1375_), .B(_1374_), .S(_2463_), .Y(_1376_) );
	NOR2X1 NOR2X1_123 ( .A(_1373__bF_buf3), .B(_1376_), .Y(_1377_) );
	OAI21X1 OAI21X1_372 ( .A(concatenador_count_1_bF_buf2), .B(concatenador_count_2_), .C(concatenador_count_3_), .Y(_1378_) );
	OAI21X1 OAI21X1_373 ( .A(_2465_), .B(concatenador_count_1_bF_buf1), .C(_1378_), .Y(_1379_) );
	XNOR2X1 XNOR2X1_24 ( .A(concatenador_count_1_bF_buf0), .B(concatenador_count_2_), .Y(_1380_) );
	MUX2X1 MUX2X1_4 ( .A(micro_hash_synth_W_25__0_), .B(micro_hash_synth_W_24__0_), .S(concatenador_count_0_bF_buf5), .Y(_1381_) );
	MUX2X1 MUX2X1_5 ( .A(micro_hash_synth_W_27__0_), .B(micro_hash_synth_W_26__0_), .S(concatenador_count_0_bF_buf4), .Y(_1382_) );
	MUX2X1 MUX2X1_6 ( .A(_1382_), .B(_1381_), .S(_2463_), .Y(_1383_) );
	OAI21X1 OAI21X1_374 ( .A(_1383_), .B(_1380__bF_buf6), .C(_1379__bF_buf3), .Y(_1384_) );
	MUX2X1 MUX2X1_7 ( .A(micro_hash_synth_W_23__0_), .B(micro_hash_synth_W_22__0_), .S(concatenador_count_0_bF_buf3), .Y(_1385_) );
	MUX2X1 MUX2X1_8 ( .A(micro_hash_synth_W_21__0_), .B(micro_hash_synth_W_20__0_), .S(concatenador_count_0_bF_buf2), .Y(_1386_) );
	MUX2X1 MUX2X1_9 ( .A(_1386_), .B(_1385_), .S(concatenador_count_1_bF_buf6), .Y(_1387_) );
	NOR2X1 NOR2X1_124 ( .A(_1373__bF_buf2), .B(_1387_), .Y(_1388_) );
	AND2X2 AND2X2_34 ( .A(_1370_), .B(_1378_), .Y(_1389_) );
	MUX2X1 MUX2X1_10 ( .A(micro_hash_synth_W_19__0_), .B(micro_hash_synth_W_18__0_), .S(concatenador_count_0_bF_buf1), .Y(_1390_) );
	MUX2X1 MUX2X1_11 ( .A(micro_hash_synth_W_17__0_), .B(micro_hash_synth_W_16__0_), .S(concatenador_count_0_bF_buf0), .Y(_1391_) );
	MUX2X1 MUX2X1_12 ( .A(_1391_), .B(_1390_), .S(concatenador_count_1_bF_buf5), .Y(_1392_) );
	OAI21X1 OAI21X1_375 ( .A(_1392_), .B(_1380__bF_buf5), .C(_1389_), .Y(_1393_) );
	OAI22X1 OAI22X1_56 ( .A(_1384_), .B(_1377_), .C(_1388_), .D(_1393_), .Y(_1394_) );
	MUX2X1 MUX2X1_13 ( .A(micro_hash_synth_W_15__0_), .B(micro_hash_synth_W_14__0_), .S(concatenador_count_0_bF_buf11), .Y(_1395_) );
	MUX2X1 MUX2X1_14 ( .A(micro_hash_synth_W_13__0_), .B(micro_hash_synth_W_12__0_), .S(concatenador_count_0_bF_buf10), .Y(_1396_) );
	MUX2X1 MUX2X1_15 ( .A(_1396_), .B(_1395_), .S(concatenador_count_1_bF_buf4), .Y(_1397_) );
	NOR2X1 NOR2X1_125 ( .A(_1373__bF_buf1), .B(_1397_), .Y(_1398_) );
	MUX2X1 MUX2X1_16 ( .A(micro_hash_synth_W_11__0_), .B(micro_hash_synth_W_10__0_), .S(concatenador_count_0_bF_buf9), .Y(_1399_) );
	MUX2X1 MUX2X1_17 ( .A(micro_hash_synth_W_9__0_), .B(micro_hash_synth_W_8__0_), .S(concatenador_count_0_bF_buf8), .Y(_1400_) );
	MUX2X1 MUX2X1_18 ( .A(_1400_), .B(_1399_), .S(concatenador_count_1_bF_buf3), .Y(_1401_) );
	OAI21X1 OAI21X1_376 ( .A(_1401_), .B(_1380__bF_buf4), .C(_1379__bF_buf2), .Y(_1402_) );
	MUX2X1 MUX2X1_19 ( .A(micro_hash_synth_W_7__0_), .B(micro_hash_synth_W_6__0_), .S(concatenador_count_0_bF_buf7), .Y(_1403_) );
	MUX2X1 MUX2X1_20 ( .A(micro_hash_synth_W_5__0_), .B(micro_hash_synth_W_4__0_), .S(concatenador_count_0_bF_buf6), .Y(_1404_) );
	MUX2X1 MUX2X1_21 ( .A(_1404_), .B(_1403_), .S(concatenador_count_1_bF_buf2), .Y(_1405_) );
	NOR2X1 NOR2X1_126 ( .A(_1373__bF_buf0), .B(_1405_), .Y(_1406_) );
	MUX2X1 MUX2X1_22 ( .A(micro_hash_synth_W_3__0_), .B(micro_hash_synth_W_2__0_), .S(concatenador_count_0_bF_buf5), .Y(_1407_) );
	MUX2X1 MUX2X1_23 ( .A(micro_hash_synth_W_1__0_), .B(micro_hash_synth_W_0__0_), .S(concatenador_count_0_bF_buf4), .Y(_1408_) );
	MUX2X1 MUX2X1_24 ( .A(_1408_), .B(_1407_), .S(concatenador_count_1_bF_buf1), .Y(_1409_) );
	OAI21X1 OAI21X1_377 ( .A(_1409_), .B(_1380__bF_buf3), .C(_1389_), .Y(_1410_) );
	OAI22X1 OAI22X1_57 ( .A(_1402_), .B(_1398_), .C(_1406_), .D(_1410_), .Y(_1411_) );
	MUX2X1 MUX2X1_25 ( .A(_1411_), .B(_1394_), .S(_1372_), .Y(_1412_) );
	NOR2X1 NOR2X1_127 ( .A(_1369_), .B(_1412_), .Y(_1413_) );
	INVX1 INVX1_371 ( .A(_1412_), .Y(_1414_) );
	NOR2X1 NOR2X1_128 ( .A(_1205__bF_buf2), .B(_1366_), .Y(_1415_) );
	OAI21X1 OAI21X1_378 ( .A(_1414_), .B(_1368_), .C(_1415_), .Y(_1416_) );
	OAI22X1 OAI22X1_58 ( .A(_1367_), .B(_1356_), .C(_1416_), .D(_1413_), .Y(_930__0_) );
	NAND2X1 NAND2X1_134 ( .A(micro_hash_synth_k_0_), .B(micro_hash_synth_x_0_), .Y(_1417_) );
	OAI21X1 OAI21X1_379 ( .A(_1412_), .B(_1369_), .C(_1417_), .Y(_1418_) );
	INVX1 INVX1_372 ( .A(micro_hash_synth_x_1_), .Y(_1419_) );
	NOR2X1 NOR2X1_129 ( .A(_1357_), .B(_1419_), .Y(_1420_) );
	NOR2X1 NOR2X1_130 ( .A(micro_hash_synth_k_1_), .B(micro_hash_synth_x_1_), .Y(_1421_) );
	NAND2X1 NAND2X1_135 ( .A(concatenador_count_0_bF_buf3), .B(micro_hash_synth_W_23__1_), .Y(_1422_) );
	OAI21X1 OAI21X1_380 ( .A(_2576_), .B(concatenador_count_0_bF_buf2), .C(_1422_), .Y(_1423_) );
	INVX1 INVX1_373 ( .A(micro_hash_synth_W_20__1_), .Y(_1424_) );
	NAND2X1 NAND2X1_136 ( .A(concatenador_count_0_bF_buf1), .B(micro_hash_synth_W_21__1_), .Y(_1425_) );
	OAI21X1 OAI21X1_381 ( .A(_1424_), .B(concatenador_count_0_bF_buf0), .C(_1425_), .Y(_1426_) );
	MUX2X1 MUX2X1_26 ( .A(_1426_), .B(_1423_), .S(concatenador_count_1_bF_buf0), .Y(_1427_) );
	AND2X2 AND2X2_35 ( .A(_1427_), .B(_1380__bF_buf2), .Y(_1428_) );
	INVX1 INVX1_374 ( .A(micro_hash_synth_W_16__1_), .Y(_1429_) );
	NAND2X1 NAND2X1_137 ( .A(concatenador_count_1_bF_buf6), .B(_2462_), .Y(_1430_) );
	OAI21X1 OAI21X1_382 ( .A(_1429_), .B(_1430_), .C(_1373__bF_buf3), .Y(_1431_) );
	INVX1 INVX1_375 ( .A(micro_hash_synth_W_17__1_), .Y(_1432_) );
	NAND2X1 NAND2X1_138 ( .A(concatenador_count_0_bF_buf11), .B(concatenador_count_1_bF_buf5), .Y(_1433_) );
	MUX2X1 MUX2X1_27 ( .A(micro_hash_synth_W_19__1_), .B(micro_hash_synth_W_18__1_), .S(concatenador_count_0_bF_buf10), .Y(_1434_) );
	OAI22X1 OAI22X1_59 ( .A(_1432_), .B(_1433_), .C(_1434_), .D(concatenador_count_1_bF_buf4), .Y(_1435_) );
	OAI21X1 OAI21X1_383 ( .A(_1431_), .B(_1435_), .C(_1389_), .Y(_1436_) );
	NOR2X1 NOR2X1_131 ( .A(_1436_), .B(_1428_), .Y(_1437_) );
	INVX1 INVX1_376 ( .A(micro_hash_synth_W_28__1_), .Y(_1438_) );
	NAND2X1 NAND2X1_139 ( .A(concatenador_count_0_bF_buf9), .B(micro_hash_synth_W_29__1_), .Y(_1439_) );
	OAI21X1 OAI21X1_384 ( .A(_1438_), .B(concatenador_count_0_bF_buf8), .C(_1439_), .Y(_1440_) );
	INVX1 INVX1_377 ( .A(micro_hash_synth_W_30__1_), .Y(_1441_) );
	NAND2X1 NAND2X1_140 ( .A(concatenador_count_0_bF_buf7), .B(micro_hash_synth_W_31__1_), .Y(_1442_) );
	OAI21X1 OAI21X1_385 ( .A(_1441_), .B(concatenador_count_0_bF_buf6), .C(_1442_), .Y(_1443_) );
	MUX2X1 MUX2X1_28 ( .A(_1443_), .B(_1440_), .S(_2463_), .Y(_1444_) );
	AND2X2 AND2X2_36 ( .A(_1444_), .B(_1380__bF_buf1), .Y(_1445_) );
	MUX2X1 MUX2X1_29 ( .A(micro_hash_synth_W_25__1_), .B(micro_hash_synth_W_24__1_), .S(concatenador_count_0_bF_buf5), .Y(_1446_) );
	MUX2X1 MUX2X1_30 ( .A(micro_hash_synth_W_27__1_), .B(micro_hash_synth_W_26__1_), .S(concatenador_count_0_bF_buf4), .Y(_1447_) );
	MUX2X1 MUX2X1_31 ( .A(_1447_), .B(_1446_), .S(_2463_), .Y(_1448_) );
	OAI21X1 OAI21X1_386 ( .A(_1448_), .B(_1380__bF_buf0), .C(_1379__bF_buf1), .Y(_1449_) );
	OAI21X1 OAI21X1_387 ( .A(_1445_), .B(_1449_), .C(_1371_), .Y(_1450_) );
	INVX1 INVX1_378 ( .A(micro_hash_synth_W_4__1_), .Y(_1451_) );
	OAI21X1 OAI21X1_388 ( .A(_1451_), .B(_1430_), .C(_1380__bF_buf6), .Y(_1452_) );
	INVX1 INVX1_379 ( .A(micro_hash_synth_W_5__1_), .Y(_1453_) );
	MUX2X1 MUX2X1_32 ( .A(micro_hash_synth_W_7__1_), .B(micro_hash_synth_W_6__1_), .S(concatenador_count_0_bF_buf3), .Y(_1454_) );
	OAI22X1 OAI22X1_60 ( .A(_1453_), .B(_1433_), .C(_1454_), .D(concatenador_count_1_bF_buf3), .Y(_1455_) );
	MUX2X1 MUX2X1_33 ( .A(micro_hash_synth_W_1__1_), .B(micro_hash_synth_W_0__1_), .S(concatenador_count_0_bF_buf2), .Y(_1456_) );
	MUX2X1 MUX2X1_34 ( .A(micro_hash_synth_W_3__1_), .B(micro_hash_synth_W_2__1_), .S(concatenador_count_0_bF_buf1), .Y(_1457_) );
	MUX2X1 MUX2X1_35 ( .A(_1457_), .B(_1456_), .S(_2463_), .Y(_1458_) );
	OAI22X1 OAI22X1_61 ( .A(_1380__bF_buf5), .B(_1458_), .C(_1452_), .D(_1455_), .Y(_1459_) );
	OAI21X1 OAI21X1_389 ( .A(_2535_), .B(_1430_), .C(_1380__bF_buf4), .Y(_1460_) );
	MUX2X1 MUX2X1_36 ( .A(micro_hash_synth_W_15__1_), .B(micro_hash_synth_W_14__1_), .S(concatenador_count_0_bF_buf0), .Y(_1461_) );
	OAI22X1 OAI22X1_62 ( .A(_2479_), .B(_1433_), .C(_1461_), .D(concatenador_count_1_bF_buf2), .Y(_1462_) );
	NOR2X1 NOR2X1_132 ( .A(_1462_), .B(_1460_), .Y(_1463_) );
	INVX1 INVX1_380 ( .A(micro_hash_synth_W_8__1_), .Y(_1464_) );
	OAI21X1 OAI21X1_390 ( .A(_1464_), .B(_1430_), .C(_1373__bF_buf2), .Y(_1465_) );
	MUX2X1 MUX2X1_37 ( .A(micro_hash_synth_W_11__1_), .B(micro_hash_synth_W_10__1_), .S(concatenador_count_0_bF_buf11), .Y(_1466_) );
	OAI22X1 OAI22X1_63 ( .A(_2515_), .B(_1433_), .C(_1466_), .D(concatenador_count_1_bF_buf1), .Y(_1467_) );
	OAI21X1 OAI21X1_391 ( .A(_1465_), .B(_1467_), .C(_1379__bF_buf0), .Y(_1468_) );
	OAI22X1 OAI22X1_64 ( .A(_1468_), .B(_1463_), .C(_1459_), .D(_1379__bF_buf3), .Y(_1469_) );
	OAI22X1 OAI22X1_65 ( .A(_1450_), .B(_1437_), .C(_1371_), .D(_1469_), .Y(_1470_) );
	OAI21X1 OAI21X1_392 ( .A(_1420_), .B(_1421_), .C(_1470_), .Y(_1471_) );
	NOR2X1 NOR2X1_133 ( .A(_1421_), .B(_1420_), .Y(_1472_) );
	INVX1 INVX1_381 ( .A(micro_hash_synth_W_18__1_), .Y(_1473_) );
	NAND2X1 NAND2X1_141 ( .A(concatenador_count_0_bF_buf10), .B(micro_hash_synth_W_19__1_), .Y(_1474_) );
	OAI21X1 OAI21X1_393 ( .A(_1473_), .B(concatenador_count_0_bF_buf9), .C(_1474_), .Y(_1475_) );
	NAND2X1 NAND2X1_142 ( .A(concatenador_count_0_bF_buf8), .B(micro_hash_synth_W_17__1_), .Y(_1476_) );
	OAI21X1 OAI21X1_394 ( .A(_1429_), .B(concatenador_count_0_bF_buf7), .C(_1476_), .Y(_1477_) );
	MUX2X1 MUX2X1_38 ( .A(_1477_), .B(_1475_), .S(concatenador_count_1_bF_buf0), .Y(_1478_) );
	MUX2X1 MUX2X1_39 ( .A(_1427_), .B(_1478_), .S(_1380__bF_buf3), .Y(_1479_) );
	NAND2X1 NAND2X1_143 ( .A(concatenador_count_0_bF_buf6), .B(micro_hash_synth_W_25__1_), .Y(_1480_) );
	OAI21X1 OAI21X1_395 ( .A(_2480_), .B(concatenador_count_0_bF_buf5), .C(_1480_), .Y(_1481_) );
	NAND2X1 NAND2X1_144 ( .A(concatenador_count_0_bF_buf4), .B(micro_hash_synth_W_27__1_), .Y(_1482_) );
	OAI21X1 OAI21X1_396 ( .A(_2534_), .B(concatenador_count_0_bF_buf3), .C(_1482_), .Y(_1483_) );
	MUX2X1 MUX2X1_40 ( .A(_1483_), .B(_1481_), .S(_2463_), .Y(_1484_) );
	MUX2X1 MUX2X1_41 ( .A(_1444_), .B(_1484_), .S(_1380__bF_buf2), .Y(_1485_) );
	MUX2X1 MUX2X1_42 ( .A(_1485_), .B(_1479_), .S(_1379__bF_buf2), .Y(_1486_) );
	INVX1 INVX1_382 ( .A(micro_hash_synth_W_6__1_), .Y(_1487_) );
	NAND2X1 NAND2X1_145 ( .A(concatenador_count_0_bF_buf2), .B(micro_hash_synth_W_7__1_), .Y(_1488_) );
	OAI21X1 OAI21X1_397 ( .A(_1487_), .B(concatenador_count_0_bF_buf1), .C(_1488_), .Y(_1489_) );
	NAND2X1 NAND2X1_146 ( .A(concatenador_count_0_bF_buf0), .B(micro_hash_synth_W_5__1_), .Y(_1490_) );
	OAI21X1 OAI21X1_398 ( .A(_1451_), .B(concatenador_count_0_bF_buf11), .C(_1490_), .Y(_1491_) );
	MUX2X1 MUX2X1_43 ( .A(_1491_), .B(_1489_), .S(concatenador_count_1_bF_buf6), .Y(_1492_) );
	INVX1 INVX1_383 ( .A(micro_hash_synth_W_0__1_), .Y(_1493_) );
	NAND2X1 NAND2X1_147 ( .A(concatenador_count_0_bF_buf10), .B(micro_hash_synth_W_1__1_), .Y(_1494_) );
	OAI21X1 OAI21X1_399 ( .A(_1493_), .B(concatenador_count_0_bF_buf9), .C(_1494_), .Y(_1495_) );
	INVX1 INVX1_384 ( .A(micro_hash_synth_W_2__1_), .Y(_1496_) );
	NAND2X1 NAND2X1_148 ( .A(concatenador_count_0_bF_buf8), .B(micro_hash_synth_W_3__1_), .Y(_1497_) );
	OAI21X1 OAI21X1_400 ( .A(_1496_), .B(concatenador_count_0_bF_buf7), .C(_1497_), .Y(_1498_) );
	MUX2X1 MUX2X1_44 ( .A(_1498_), .B(_1495_), .S(_2463_), .Y(_1499_) );
	MUX2X1 MUX2X1_45 ( .A(_1492_), .B(_1499_), .S(_1380__bF_buf1), .Y(_1500_) );
	INVX1 INVX1_385 ( .A(micro_hash_synth_W_14__1_), .Y(_1501_) );
	NAND2X1 NAND2X1_149 ( .A(concatenador_count_0_bF_buf6), .B(micro_hash_synth_W_15__1_), .Y(_1502_) );
	OAI21X1 OAI21X1_401 ( .A(_1501_), .B(concatenador_count_0_bF_buf5), .C(_1502_), .Y(_1503_) );
	NAND2X1 NAND2X1_150 ( .A(concatenador_count_0_bF_buf4), .B(micro_hash_synth_W_13__1_), .Y(_1504_) );
	OAI21X1 OAI21X1_402 ( .A(_2535_), .B(concatenador_count_0_bF_buf3), .C(_1504_), .Y(_1505_) );
	MUX2X1 MUX2X1_46 ( .A(_1505_), .B(_1503_), .S(concatenador_count_1_bF_buf5), .Y(_1506_) );
	INVX1 INVX1_386 ( .A(micro_hash_synth_W_10__1_), .Y(_1507_) );
	NAND2X1 NAND2X1_151 ( .A(concatenador_count_0_bF_buf2), .B(micro_hash_synth_W_11__1_), .Y(_1508_) );
	OAI21X1 OAI21X1_403 ( .A(_1507_), .B(concatenador_count_0_bF_buf1), .C(_1508_), .Y(_1509_) );
	NAND2X1 NAND2X1_152 ( .A(concatenador_count_0_bF_buf0), .B(micro_hash_synth_W_9__1_), .Y(_1510_) );
	OAI21X1 OAI21X1_404 ( .A(_1464_), .B(concatenador_count_0_bF_buf11), .C(_1510_), .Y(_1511_) );
	MUX2X1 MUX2X1_47 ( .A(_1511_), .B(_1509_), .S(concatenador_count_1_bF_buf4), .Y(_1512_) );
	MUX2X1 MUX2X1_48 ( .A(_1506_), .B(_1512_), .S(_1380__bF_buf0), .Y(_1513_) );
	MUX2X1 MUX2X1_49 ( .A(_1513_), .B(_1500_), .S(_1379__bF_buf1), .Y(_1514_) );
	MUX2X1 MUX2X1_50 ( .A(_1514_), .B(_1486_), .S(_1372_), .Y(_1515_) );
	NAND2X1 NAND2X1_153 ( .A(_1472_), .B(_1515_), .Y(_1516_) );
	AOI21X1 AOI21X1_304 ( .A(_1516_), .B(_1471_), .C(_1418_), .Y(_1517_) );
	NOR2X1 NOR2X1_134 ( .A(_2468_), .B(_1366_), .Y(_1518_) );
	NAND3X1 NAND3X1_76 ( .A(_1516_), .B(_1471_), .C(_1418_), .Y(_1519_) );
	NAND2X1 NAND2X1_154 ( .A(_1518_), .B(_1519_), .Y(_1520_) );
	AOI21X1 AOI21X1_305 ( .A(micro_hash_synth_c_1_), .B(_1366_), .C(_1205__bF_buf1), .Y(_1521_) );
	OAI21X1 OAI21X1_405 ( .A(_1520_), .B(_1517_), .C(_1521_), .Y(_930__1_) );
	INVX1 INVX1_387 ( .A(_1518_), .Y(_1522_) );
	INVX1 INVX1_388 ( .A(_1420_), .Y(_1523_) );
	OAI21X1 OAI21X1_406 ( .A(_1470_), .B(_1421_), .C(_1523_), .Y(_1524_) );
	XOR2X1 XOR2X1_27 ( .A(micro_hash_synth_k_2_), .B(micro_hash_synth_x_2_), .Y(_1525_) );
	INVX1 INVX1_389 ( .A(_1525_), .Y(_1526_) );
	INVX1 INVX1_390 ( .A(micro_hash_synth_W_16__2_), .Y(_1527_) );
	OAI21X1 OAI21X1_407 ( .A(_1527_), .B(_1430_), .C(_1373__bF_buf1), .Y(_1528_) );
	INVX1 INVX1_391 ( .A(micro_hash_synth_W_17__2_), .Y(_1529_) );
	MUX2X1 MUX2X1_51 ( .A(micro_hash_synth_W_19__2_), .B(micro_hash_synth_W_18__2_), .S(concatenador_count_0_bF_buf10), .Y(_1530_) );
	OAI22X1 OAI22X1_66 ( .A(_1529_), .B(_1433_), .C(_1530_), .D(concatenador_count_1_bF_buf3), .Y(_1531_) );
	NOR2X1 NOR2X1_135 ( .A(_1528_), .B(_1531_), .Y(_1532_) );
	MUX2X1 MUX2X1_52 ( .A(micro_hash_synth_W_23__2_), .B(micro_hash_synth_W_22__2_), .S(concatenador_count_0_bF_buf9), .Y(_1533_) );
	MUX2X1 MUX2X1_53 ( .A(micro_hash_synth_W_21__2_), .B(micro_hash_synth_W_20__2_), .S(concatenador_count_0_bF_buf8), .Y(_1534_) );
	MUX2X1 MUX2X1_54 ( .A(_1534_), .B(_1533_), .S(concatenador_count_1_bF_buf2), .Y(_1535_) );
	OAI21X1 OAI21X1_408 ( .A(_1535_), .B(_1373__bF_buf0), .C(_1389_), .Y(_1536_) );
	NOR2X1 NOR2X1_136 ( .A(_1536_), .B(_1532_), .Y(_1537_) );
	MUX2X1 MUX2X1_55 ( .A(micro_hash_synth_W_29__2_), .B(micro_hash_synth_W_28__2_), .S(concatenador_count_0_bF_buf7), .Y(_1538_) );
	MUX2X1 MUX2X1_56 ( .A(micro_hash_synth_W_31__2_), .B(micro_hash_synth_W_30__2_), .S(concatenador_count_0_bF_buf6), .Y(_1539_) );
	MUX2X1 MUX2X1_57 ( .A(_1539_), .B(_1538_), .S(_2463_), .Y(_1540_) );
	NOR2X1 NOR2X1_137 ( .A(_1373__bF_buf3), .B(_1540_), .Y(_1541_) );
	MUX2X1 MUX2X1_58 ( .A(micro_hash_synth_W_25__2_), .B(micro_hash_synth_W_24__2_), .S(concatenador_count_0_bF_buf5), .Y(_1542_) );
	MUX2X1 MUX2X1_59 ( .A(micro_hash_synth_W_27__2_), .B(micro_hash_synth_W_26__2_), .S(concatenador_count_0_bF_buf4), .Y(_1543_) );
	MUX2X1 MUX2X1_60 ( .A(_1543_), .B(_1542_), .S(_2463_), .Y(_1544_) );
	OAI21X1 OAI21X1_409 ( .A(_1544_), .B(_1380__bF_buf6), .C(_1379__bF_buf0), .Y(_1545_) );
	OAI21X1 OAI21X1_410 ( .A(_1545_), .B(_1541_), .C(_1371_), .Y(_1546_) );
	INVX4 INVX4_9 ( .A(_1433_), .Y(_1547_) );
	AOI22X1 AOI22X1_28 ( .A(micro_hash_synth_W_13__2_), .B(_1547__bF_buf3), .C(_2609__bF_buf2), .D(micro_hash_synth_W_12__2_), .Y(_1548_) );
	NOR2X1 NOR2X1_138 ( .A(concatenador_count_1_bF_buf1), .B(_2462_), .Y(_1549_) );
	AOI22X1 AOI22X1_29 ( .A(micro_hash_synth_W_14__2_), .B(_2470__bF_buf0), .C(_1549__bF_buf3), .D(micro_hash_synth_W_15__2_), .Y(_1550_) );
	AND2X2 AND2X2_37 ( .A(_1548_), .B(_1550_), .Y(_1551_) );
	MUX2X1 MUX2X1_61 ( .A(micro_hash_synth_W_11__2_), .B(micro_hash_synth_W_10__2_), .S(concatenador_count_0_bF_buf3), .Y(_1552_) );
	MUX2X1 MUX2X1_62 ( .A(micro_hash_synth_W_9__2_), .B(micro_hash_synth_W_8__2_), .S(concatenador_count_0_bF_buf2), .Y(_1553_) );
	MUX2X1 MUX2X1_63 ( .A(_1553_), .B(_1552_), .S(concatenador_count_1_bF_buf0), .Y(_1554_) );
	OAI21X1 OAI21X1_411 ( .A(_1554_), .B(_1380__bF_buf5), .C(_1379__bF_buf3), .Y(_1555_) );
	AOI21X1 AOI21X1_306 ( .A(_1380__bF_buf4), .B(_1551_), .C(_1555_), .Y(_1556_) );
	INVX1 INVX1_392 ( .A(micro_hash_synth_W_6__2_), .Y(_1557_) );
	NAND2X1 NAND2X1_155 ( .A(concatenador_count_0_bF_buf1), .B(micro_hash_synth_W_7__2_), .Y(_1558_) );
	OAI21X1 OAI21X1_412 ( .A(_1557_), .B(concatenador_count_0_bF_buf0), .C(_1558_), .Y(_1559_) );
	INVX1 INVX1_393 ( .A(micro_hash_synth_W_4__2_), .Y(_1560_) );
	NAND2X1 NAND2X1_156 ( .A(concatenador_count_0_bF_buf11), .B(micro_hash_synth_W_5__2_), .Y(_1561_) );
	OAI21X1 OAI21X1_413 ( .A(_1560_), .B(concatenador_count_0_bF_buf10), .C(_1561_), .Y(_1562_) );
	MUX2X1 MUX2X1_64 ( .A(_1562_), .B(_1559_), .S(concatenador_count_1_bF_buf6), .Y(_1563_) );
	AND2X2 AND2X2_38 ( .A(_1563_), .B(_1380__bF_buf3), .Y(_1564_) );
	MUX2X1 MUX2X1_65 ( .A(micro_hash_synth_W_3__2_), .B(micro_hash_synth_W_2__2_), .S(concatenador_count_0_bF_buf9), .Y(_1565_) );
	MUX2X1 MUX2X1_66 ( .A(micro_hash_synth_W_1__2_), .B(micro_hash_synth_W_0__2_), .S(concatenador_count_0_bF_buf8), .Y(_1566_) );
	MUX2X1 MUX2X1_67 ( .A(_1566_), .B(_1565_), .S(concatenador_count_1_bF_buf5), .Y(_1567_) );
	OAI21X1 OAI21X1_414 ( .A(_1567_), .B(_1380__bF_buf2), .C(_1389_), .Y(_1568_) );
	OAI21X1 OAI21X1_415 ( .A(_1564_), .B(_1568_), .C(_1372_), .Y(_1569_) );
	OAI22X1 OAI22X1_67 ( .A(_1537_), .B(_1546_), .C(_1569_), .D(_1556_), .Y(_1570_) );
	NAND2X1 NAND2X1_157 ( .A(_1526_), .B(_1570_), .Y(_1571_) );
	OR2X2 OR2X2_26 ( .A(_1546_), .B(_1537_), .Y(_1572_) );
	NAND3X1 NAND3X1_77 ( .A(_1380__bF_buf1), .B(_1550_), .C(_1548_), .Y(_1573_) );
	OR2X2 OR2X2_27 ( .A(_1554_), .B(_1380__bF_buf0), .Y(_1574_) );
	NAND3X1 NAND3X1_78 ( .A(_1379__bF_buf2), .B(_1573_), .C(_1574_), .Y(_1575_) );
	AND2X2 AND2X2_39 ( .A(_1567_), .B(_1373__bF_buf2), .Y(_1576_) );
	NOR2X1 NOR2X1_139 ( .A(_1373__bF_buf1), .B(_1563_), .Y(_1577_) );
	OAI21X1 OAI21X1_416 ( .A(_1577_), .B(_1576_), .C(_1389_), .Y(_1578_) );
	NAND3X1 NAND3X1_79 ( .A(_1372_), .B(_1575_), .C(_1578_), .Y(_1579_) );
	NAND3X1 NAND3X1_80 ( .A(_1525_), .B(_1579_), .C(_1572_), .Y(_1580_) );
	NAND3X1 NAND3X1_81 ( .A(_1571_), .B(_1580_), .C(_1524_), .Y(_1581_) );
	AOI21X1 AOI21X1_307 ( .A(_1472_), .B(_1515_), .C(_1420_), .Y(_1582_) );
	AOI21X1 AOI21X1_308 ( .A(_1579_), .B(_1572_), .C(_1525_), .Y(_1583_) );
	NOR2X1 NOR2X1_140 ( .A(_1526_), .B(_1570_), .Y(_1584_) );
	OAI21X1 OAI21X1_417 ( .A(_1583_), .B(_1584_), .C(_1582_), .Y(_1585_) );
	NAND2X1 NAND2X1_158 ( .A(_1585_), .B(_1581_), .Y(_1586_) );
	NAND2X1 NAND2X1_159 ( .A(_1519_), .B(_1586_), .Y(_1587_) );
	OAI21X1 OAI21X1_418 ( .A(_1583_), .B(_1584_), .C(_1524_), .Y(_1588_) );
	NAND3X1 NAND3X1_82 ( .A(_1571_), .B(_1580_), .C(_1582_), .Y(_1589_) );
	AOI21X1 AOI21X1_309 ( .A(_1588_), .B(_1589_), .C(_1519_), .Y(_1590_) );
	INVX1 INVX1_394 ( .A(_1590_), .Y(_1591_) );
	NAND2X1 NAND2X1_160 ( .A(_1587_), .B(_1591_), .Y(_1592_) );
	AOI21X1 AOI21X1_310 ( .A(micro_hash_synth_c_2_), .B(_1366_), .C(_1205__bF_buf0), .Y(_1593_) );
	OAI21X1 OAI21X1_419 ( .A(_1592_), .B(_1522_), .C(_1593_), .Y(_930__2_) );
	OAI21X1 OAI21X1_420 ( .A(_1586_), .B(_1519_), .C(_1581_), .Y(_1594_) );
	INVX1 INVX1_395 ( .A(micro_hash_synth_x_2_), .Y(_1595_) );
	OAI21X1 OAI21X1_421 ( .A(_1358_), .B(_1595_), .C(_1580_), .Y(_1596_) );
	NOR2X1 NOR2X1_141 ( .A(micro_hash_synth_k_3_), .B(micro_hash_synth_x_3_), .Y(_1597_) );
	NAND2X1 NAND2X1_161 ( .A(micro_hash_synth_k_3_), .B(micro_hash_synth_x_3_), .Y(_1598_) );
	INVX1 INVX1_396 ( .A(_1598_), .Y(_1599_) );
	NOR2X1 NOR2X1_142 ( .A(_1597_), .B(_1599_), .Y(_1600_) );
	NAND2X1 NAND2X1_162 ( .A(concatenador_count_0_bF_buf7), .B(micro_hash_synth_W_23__3_), .Y(_1601_) );
	OAI21X1 OAI21X1_422 ( .A(_2586_), .B(concatenador_count_0_bF_buf6), .C(_1601_), .Y(_1602_) );
	INVX1 INVX1_397 ( .A(micro_hash_synth_W_20__3_), .Y(_1603_) );
	NAND2X1 NAND2X1_163 ( .A(concatenador_count_0_bF_buf5), .B(micro_hash_synth_W_21__3_), .Y(_1604_) );
	OAI21X1 OAI21X1_423 ( .A(_1603_), .B(concatenador_count_0_bF_buf4), .C(_1604_), .Y(_1605_) );
	MUX2X1 MUX2X1_68 ( .A(_1605_), .B(_1602_), .S(concatenador_count_1_bF_buf4), .Y(_1606_) );
	INVX1 INVX1_398 ( .A(micro_hash_synth_W_18__3_), .Y(_1607_) );
	NAND2X1 NAND2X1_164 ( .A(concatenador_count_0_bF_buf3), .B(micro_hash_synth_W_19__3_), .Y(_1608_) );
	OAI21X1 OAI21X1_424 ( .A(_1607_), .B(concatenador_count_0_bF_buf2), .C(_1608_), .Y(_1609_) );
	INVX1 INVX1_399 ( .A(micro_hash_synth_W_16__3_), .Y(_1610_) );
	NAND2X1 NAND2X1_165 ( .A(concatenador_count_0_bF_buf1), .B(micro_hash_synth_W_17__3_), .Y(_1611_) );
	OAI21X1 OAI21X1_425 ( .A(_1610_), .B(concatenador_count_0_bF_buf0), .C(_1611_), .Y(_1612_) );
	MUX2X1 MUX2X1_69 ( .A(_1612_), .B(_1609_), .S(concatenador_count_1_bF_buf3), .Y(_1613_) );
	MUX2X1 MUX2X1_70 ( .A(_1606_), .B(_1613_), .S(_1380__bF_buf6), .Y(_1614_) );
	INVX1 INVX1_400 ( .A(micro_hash_synth_W_30__3_), .Y(_1615_) );
	NAND2X1 NAND2X1_166 ( .A(concatenador_count_0_bF_buf11), .B(micro_hash_synth_W_31__3_), .Y(_1616_) );
	OAI21X1 OAI21X1_426 ( .A(_1615_), .B(concatenador_count_0_bF_buf10), .C(_1616_), .Y(_1617_) );
	INVX1 INVX1_401 ( .A(micro_hash_synth_W_28__3_), .Y(_1618_) );
	NAND2X1 NAND2X1_167 ( .A(concatenador_count_0_bF_buf9), .B(micro_hash_synth_W_29__3_), .Y(_1619_) );
	OAI21X1 OAI21X1_427 ( .A(_1618_), .B(concatenador_count_0_bF_buf8), .C(_1619_), .Y(_1620_) );
	MUX2X1 MUX2X1_71 ( .A(_1620_), .B(_1617_), .S(concatenador_count_1_bF_buf2), .Y(_1621_) );
	NAND2X1 NAND2X1_168 ( .A(concatenador_count_0_bF_buf7), .B(micro_hash_synth_W_27__3_), .Y(_1622_) );
	OAI21X1 OAI21X1_428 ( .A(_2544_), .B(concatenador_count_0_bF_buf6), .C(_1622_), .Y(_1623_) );
	NAND2X1 NAND2X1_169 ( .A(concatenador_count_0_bF_buf5), .B(micro_hash_synth_W_25__3_), .Y(_1624_) );
	OAI21X1 OAI21X1_429 ( .A(_2490_), .B(concatenador_count_0_bF_buf4), .C(_1624_), .Y(_1625_) );
	MUX2X1 MUX2X1_72 ( .A(_1625_), .B(_1623_), .S(concatenador_count_1_bF_buf1), .Y(_1626_) );
	MUX2X1 MUX2X1_73 ( .A(_1621_), .B(_1626_), .S(_1380__bF_buf5), .Y(_1627_) );
	MUX2X1 MUX2X1_74 ( .A(_1627_), .B(_1614_), .S(_1379__bF_buf1), .Y(_1628_) );
	INVX1 INVX1_402 ( .A(micro_hash_synth_W_6__3_), .Y(_1629_) );
	NAND2X1 NAND2X1_170 ( .A(concatenador_count_0_bF_buf3), .B(micro_hash_synth_W_7__3_), .Y(_1630_) );
	OAI21X1 OAI21X1_430 ( .A(_1629_), .B(concatenador_count_0_bF_buf2), .C(_1630_), .Y(_1631_) );
	INVX1 INVX1_403 ( .A(micro_hash_synth_W_4__3_), .Y(_1632_) );
	NAND2X1 NAND2X1_171 ( .A(concatenador_count_0_bF_buf1), .B(micro_hash_synth_W_5__3_), .Y(_1633_) );
	OAI21X1 OAI21X1_431 ( .A(_1632_), .B(concatenador_count_0_bF_buf0), .C(_1633_), .Y(_1634_) );
	MUX2X1 MUX2X1_75 ( .A(_1634_), .B(_1631_), .S(concatenador_count_1_bF_buf0), .Y(_1635_) );
	INVX1 INVX1_404 ( .A(micro_hash_synth_W_2__3_), .Y(_1636_) );
	NAND2X1 NAND2X1_172 ( .A(concatenador_count_0_bF_buf11), .B(micro_hash_synth_W_3__3_), .Y(_1637_) );
	OAI21X1 OAI21X1_432 ( .A(_1636_), .B(concatenador_count_0_bF_buf10), .C(_1637_), .Y(_1638_) );
	INVX1 INVX1_405 ( .A(micro_hash_synth_W_0__3_), .Y(_1639_) );
	NAND2X1 NAND2X1_173 ( .A(concatenador_count_0_bF_buf9), .B(micro_hash_synth_W_1__3_), .Y(_1640_) );
	OAI21X1 OAI21X1_433 ( .A(_1639_), .B(concatenador_count_0_bF_buf8), .C(_1640_), .Y(_1641_) );
	MUX2X1 MUX2X1_76 ( .A(_1641_), .B(_1638_), .S(concatenador_count_1_bF_buf6), .Y(_1642_) );
	MUX2X1 MUX2X1_77 ( .A(_1635_), .B(_1642_), .S(_1380__bF_buf4), .Y(_1643_) );
	INVX1 INVX1_406 ( .A(micro_hash_synth_W_14__3_), .Y(_1644_) );
	NAND2X1 NAND2X1_174 ( .A(concatenador_count_0_bF_buf7), .B(micro_hash_synth_W_15__3_), .Y(_1645_) );
	OAI21X1 OAI21X1_434 ( .A(_1644_), .B(concatenador_count_0_bF_buf6), .C(_1645_), .Y(_1646_) );
	NAND2X1 NAND2X1_175 ( .A(concatenador_count_0_bF_buf5), .B(micro_hash_synth_W_13__3_), .Y(_1647_) );
	OAI21X1 OAI21X1_435 ( .A(_2545_), .B(concatenador_count_0_bF_buf4), .C(_1647_), .Y(_1648_) );
	MUX2X1 MUX2X1_78 ( .A(_1648_), .B(_1646_), .S(concatenador_count_1_bF_buf5), .Y(_1649_) );
	INVX1 INVX1_407 ( .A(micro_hash_synth_W_10__3_), .Y(_1650_) );
	NAND2X1 NAND2X1_176 ( .A(concatenador_count_0_bF_buf3), .B(micro_hash_synth_W_11__3_), .Y(_1651_) );
	OAI21X1 OAI21X1_436 ( .A(_1650_), .B(concatenador_count_0_bF_buf2), .C(_1651_), .Y(_1652_) );
	INVX1 INVX1_408 ( .A(micro_hash_synth_W_8__3_), .Y(_1653_) );
	NAND2X1 NAND2X1_177 ( .A(concatenador_count_0_bF_buf1), .B(micro_hash_synth_W_9__3_), .Y(_1654_) );
	OAI21X1 OAI21X1_437 ( .A(_1653_), .B(concatenador_count_0_bF_buf0), .C(_1654_), .Y(_1655_) );
	MUX2X1 MUX2X1_79 ( .A(_1655_), .B(_1652_), .S(concatenador_count_1_bF_buf4), .Y(_1656_) );
	MUX2X1 MUX2X1_80 ( .A(_1649_), .B(_1656_), .S(_1380__bF_buf3), .Y(_1657_) );
	MUX2X1 MUX2X1_81 ( .A(_1657_), .B(_1643_), .S(_1379__bF_buf0), .Y(_1658_) );
	MUX2X1 MUX2X1_82 ( .A(_1658_), .B(_1628_), .S(_1372_), .Y(_1659_) );
	XOR2X1 XOR2X1_28 ( .A(_1659_), .B(_1600_), .Y(_1660_) );
	NAND2X1 NAND2X1_178 ( .A(_1660_), .B(_1596_), .Y(_1661_) );
	AOI21X1 AOI21X1_311 ( .A(micro_hash_synth_k_2_), .B(micro_hash_synth_x_2_), .C(_1584_), .Y(_1662_) );
	XNOR2X1 XNOR2X1_25 ( .A(_1659_), .B(_1600_), .Y(_1663_) );
	NAND2X1 NAND2X1_179 ( .A(_1663_), .B(_1662_), .Y(_1664_) );
	NAND2X1 NAND2X1_180 ( .A(_1661_), .B(_1664_), .Y(_1665_) );
	XOR2X1 XOR2X1_29 ( .A(_1594_), .B(_1665_), .Y(_1666_) );
	AOI21X1 AOI21X1_312 ( .A(micro_hash_synth_c_3_), .B(_1366_), .C(_1205__bF_buf3), .Y(_1667_) );
	OAI21X1 OAI21X1_438 ( .A(_1666_), .B(_1522_), .C(_1667_), .Y(_930__3_) );
	AND2X2 AND2X2_40 ( .A(_1621_), .B(_1380__bF_buf2), .Y(_1668_) );
	MUX2X1 MUX2X1_83 ( .A(micro_hash_synth_W_27__3_), .B(micro_hash_synth_W_26__3_), .S(concatenador_count_0_bF_buf11), .Y(_1669_) );
	MUX2X1 MUX2X1_84 ( .A(micro_hash_synth_W_25__3_), .B(micro_hash_synth_W_24__3_), .S(concatenador_count_0_bF_buf10), .Y(_1670_) );
	MUX2X1 MUX2X1_85 ( .A(_1670_), .B(_1669_), .S(concatenador_count_1_bF_buf3), .Y(_1671_) );
	OAI21X1 OAI21X1_439 ( .A(_1671_), .B(_1380__bF_buf1), .C(_1379__bF_buf3), .Y(_1672_) );
	AND2X2 AND2X2_41 ( .A(_1606_), .B(_1380__bF_buf0), .Y(_1673_) );
	MUX2X1 MUX2X1_86 ( .A(micro_hash_synth_W_19__3_), .B(micro_hash_synth_W_18__3_), .S(concatenador_count_0_bF_buf9), .Y(_1674_) );
	MUX2X1 MUX2X1_87 ( .A(micro_hash_synth_W_17__3_), .B(micro_hash_synth_W_16__3_), .S(concatenador_count_0_bF_buf8), .Y(_1675_) );
	MUX2X1 MUX2X1_88 ( .A(_1675_), .B(_1674_), .S(concatenador_count_1_bF_buf2), .Y(_1676_) );
	OAI21X1 OAI21X1_440 ( .A(_1676_), .B(_1380__bF_buf6), .C(_1389_), .Y(_1677_) );
	OAI22X1 OAI22X1_68 ( .A(_1668_), .B(_1672_), .C(_1673_), .D(_1677_), .Y(_1678_) );
	AND2X2 AND2X2_42 ( .A(_1649_), .B(_1380__bF_buf5), .Y(_1679_) );
	MUX2X1 MUX2X1_89 ( .A(micro_hash_synth_W_11__3_), .B(micro_hash_synth_W_10__3_), .S(concatenador_count_0_bF_buf7), .Y(_1680_) );
	MUX2X1 MUX2X1_90 ( .A(micro_hash_synth_W_9__3_), .B(micro_hash_synth_W_8__3_), .S(concatenador_count_0_bF_buf6), .Y(_1681_) );
	MUX2X1 MUX2X1_91 ( .A(_1681_), .B(_1680_), .S(concatenador_count_1_bF_buf1), .Y(_1682_) );
	OAI21X1 OAI21X1_441 ( .A(_1682_), .B(_1380__bF_buf4), .C(_1379__bF_buf2), .Y(_1683_) );
	AND2X2 AND2X2_43 ( .A(_1635_), .B(_1380__bF_buf3), .Y(_1684_) );
	MUX2X1 MUX2X1_92 ( .A(micro_hash_synth_W_3__3_), .B(micro_hash_synth_W_2__3_), .S(concatenador_count_0_bF_buf5), .Y(_1685_) );
	MUX2X1 MUX2X1_93 ( .A(micro_hash_synth_W_1__3_), .B(micro_hash_synth_W_0__3_), .S(concatenador_count_0_bF_buf4), .Y(_1686_) );
	MUX2X1 MUX2X1_94 ( .A(_1686_), .B(_1685_), .S(concatenador_count_1_bF_buf0), .Y(_1687_) );
	OAI21X1 OAI21X1_442 ( .A(_1687_), .B(_1380__bF_buf2), .C(_1389_), .Y(_1688_) );
	OAI22X1 OAI22X1_69 ( .A(_1679_), .B(_1683_), .C(_1684_), .D(_1688_), .Y(_1689_) );
	MUX2X1 MUX2X1_95 ( .A(_1689_), .B(_1678_), .S(_1372_), .Y(_1690_) );
	OAI21X1 OAI21X1_443 ( .A(_1690_), .B(_1597_), .C(_1598_), .Y(_1691_) );
	INVX1 INVX1_409 ( .A(micro_hash_synth_x_4_), .Y(_1692_) );
	NAND2X1 NAND2X1_181 ( .A(_1364_), .B(_1692_), .Y(_1693_) );
	NOR2X1 NOR2X1_143 ( .A(_1364_), .B(_1692_), .Y(_1694_) );
	INVX1 INVX1_410 ( .A(_1694_), .Y(_1695_) );
	NAND2X1 NAND2X1_182 ( .A(_1693_), .B(_1695_), .Y(_1696_) );
	INVX1 INVX1_411 ( .A(micro_hash_synth_W_16__4_), .Y(_1697_) );
	NAND2X1 NAND2X1_183 ( .A(concatenador_count_0_bF_buf3), .B(micro_hash_synth_W_17__4_), .Y(_1698_) );
	OAI21X1 OAI21X1_444 ( .A(_1697_), .B(concatenador_count_0_bF_buf2), .C(_1698_), .Y(_1699_) );
	INVX1 INVX1_412 ( .A(micro_hash_synth_W_18__4_), .Y(_1700_) );
	NAND2X1 NAND2X1_184 ( .A(concatenador_count_0_bF_buf1), .B(micro_hash_synth_W_19__4_), .Y(_1701_) );
	OAI21X1 OAI21X1_445 ( .A(_1700_), .B(concatenador_count_0_bF_buf0), .C(_1701_), .Y(_1702_) );
	MUX2X1 MUX2X1_96 ( .A(_1702_), .B(_1699_), .S(_2463_), .Y(_1703_) );
	NAND2X1 NAND2X1_185 ( .A(concatenador_count_0_bF_buf11), .B(micro_hash_synth_W_23__4_), .Y(_1704_) );
	OAI21X1 OAI21X1_446 ( .A(_2591_), .B(concatenador_count_0_bF_buf10), .C(_1704_), .Y(_1705_) );
	INVX1 INVX1_413 ( .A(micro_hash_synth_W_20__4_), .Y(_1706_) );
	NAND2X1 NAND2X1_186 ( .A(concatenador_count_0_bF_buf9), .B(micro_hash_synth_W_21__4_), .Y(_1707_) );
	OAI21X1 OAI21X1_447 ( .A(_1706_), .B(concatenador_count_0_bF_buf8), .C(_1707_), .Y(_1708_) );
	MUX2X1 MUX2X1_97 ( .A(_1708_), .B(_1705_), .S(concatenador_count_1_bF_buf6), .Y(_1709_) );
	MUX2X1 MUX2X1_98 ( .A(_1709_), .B(_1703_), .S(_1380__bF_buf1), .Y(_1710_) );
	NAND2X1 NAND2X1_187 ( .A(concatenador_count_0_bF_buf7), .B(micro_hash_synth_W_27__4_), .Y(_1711_) );
	OAI21X1 OAI21X1_448 ( .A(_2549_), .B(concatenador_count_0_bF_buf6), .C(_1711_), .Y(_1712_) );
	NAND2X1 NAND2X1_188 ( .A(concatenador_count_0_bF_buf5), .B(micro_hash_synth_W_25__4_), .Y(_1713_) );
	OAI21X1 OAI21X1_449 ( .A(_2495_), .B(concatenador_count_0_bF_buf4), .C(_1713_), .Y(_1714_) );
	MUX2X1 MUX2X1_99 ( .A(_1714_), .B(_1712_), .S(concatenador_count_1_bF_buf5), .Y(_1715_) );
	INVX1 INVX1_414 ( .A(micro_hash_synth_W_30__4_), .Y(_1716_) );
	NAND2X1 NAND2X1_189 ( .A(concatenador_count_0_bF_buf3), .B(micro_hash_synth_W_31__4_), .Y(_1717_) );
	OAI21X1 OAI21X1_450 ( .A(_1716_), .B(concatenador_count_0_bF_buf2), .C(_1717_), .Y(_1718_) );
	INVX1 INVX1_415 ( .A(micro_hash_synth_W_28__4_), .Y(_1719_) );
	NAND2X1 NAND2X1_190 ( .A(concatenador_count_0_bF_buf1), .B(micro_hash_synth_W_29__4_), .Y(_1720_) );
	OAI21X1 OAI21X1_451 ( .A(_1719_), .B(concatenador_count_0_bF_buf0), .C(_1720_), .Y(_1721_) );
	MUX2X1 MUX2X1_100 ( .A(_1721_), .B(_1718_), .S(concatenador_count_1_bF_buf4), .Y(_1722_) );
	MUX2X1 MUX2X1_101 ( .A(_1722_), .B(_1715_), .S(_1380__bF_buf0), .Y(_1723_) );
	MUX2X1 MUX2X1_102 ( .A(_1723_), .B(_1710_), .S(_1379__bF_buf1), .Y(_1724_) );
	OR2X2 OR2X2_28 ( .A(_1724_), .B(_1372_), .Y(_1725_) );
	INVX1 INVX1_416 ( .A(micro_hash_synth_W_6__4_), .Y(_1726_) );
	NAND2X1 NAND2X1_191 ( .A(concatenador_count_0_bF_buf11), .B(micro_hash_synth_W_7__4_), .Y(_1727_) );
	OAI21X1 OAI21X1_452 ( .A(_1726_), .B(concatenador_count_0_bF_buf10), .C(_1727_), .Y(_1728_) );
	INVX1 INVX1_417 ( .A(micro_hash_synth_W_4__4_), .Y(_1729_) );
	NAND2X1 NAND2X1_192 ( .A(concatenador_count_0_bF_buf9), .B(micro_hash_synth_W_5__4_), .Y(_1730_) );
	OAI21X1 OAI21X1_453 ( .A(_1729_), .B(concatenador_count_0_bF_buf8), .C(_1730_), .Y(_1731_) );
	MUX2X1 MUX2X1_103 ( .A(_1731_), .B(_1728_), .S(concatenador_count_1_bF_buf3), .Y(_1732_) );
	INVX1 INVX1_418 ( .A(micro_hash_synth_W_2__4_), .Y(_1733_) );
	NAND2X1 NAND2X1_193 ( .A(concatenador_count_0_bF_buf7), .B(micro_hash_synth_W_3__4_), .Y(_1734_) );
	OAI21X1 OAI21X1_454 ( .A(_1733_), .B(concatenador_count_0_bF_buf6), .C(_1734_), .Y(_1735_) );
	INVX1 INVX1_419 ( .A(micro_hash_synth_W_0__4_), .Y(_1736_) );
	NAND2X1 NAND2X1_194 ( .A(concatenador_count_0_bF_buf5), .B(micro_hash_synth_W_1__4_), .Y(_1737_) );
	OAI21X1 OAI21X1_455 ( .A(_1736_), .B(concatenador_count_0_bF_buf4), .C(_1737_), .Y(_1738_) );
	MUX2X1 MUX2X1_104 ( .A(_1738_), .B(_1735_), .S(concatenador_count_1_bF_buf2), .Y(_1739_) );
	MUX2X1 MUX2X1_105 ( .A(_1732_), .B(_1739_), .S(_1380__bF_buf6), .Y(_1740_) );
	INVX1 INVX1_420 ( .A(micro_hash_synth_W_14__4_), .Y(_1741_) );
	NAND2X1 NAND2X1_195 ( .A(concatenador_count_0_bF_buf3), .B(micro_hash_synth_W_15__4_), .Y(_1742_) );
	OAI21X1 OAI21X1_456 ( .A(_1741_), .B(concatenador_count_0_bF_buf2), .C(_1742_), .Y(_1743_) );
	NAND2X1 NAND2X1_196 ( .A(concatenador_count_0_bF_buf1), .B(micro_hash_synth_W_13__4_), .Y(_1744_) );
	OAI21X1 OAI21X1_457 ( .A(_2550_), .B(concatenador_count_0_bF_buf0), .C(_1744_), .Y(_1745_) );
	MUX2X1 MUX2X1_106 ( .A(_1745_), .B(_1743_), .S(concatenador_count_1_bF_buf1), .Y(_1746_) );
	INVX1 INVX1_421 ( .A(micro_hash_synth_W_10__4_), .Y(_1747_) );
	NAND2X1 NAND2X1_197 ( .A(concatenador_count_0_bF_buf11), .B(micro_hash_synth_W_11__4_), .Y(_1748_) );
	OAI21X1 OAI21X1_458 ( .A(_1747_), .B(concatenador_count_0_bF_buf10), .C(_1748_), .Y(_1749_) );
	INVX1 INVX1_422 ( .A(micro_hash_synth_W_8__4_), .Y(_1750_) );
	NAND2X1 NAND2X1_198 ( .A(concatenador_count_0_bF_buf9), .B(micro_hash_synth_W_9__4_), .Y(_1751_) );
	OAI21X1 OAI21X1_459 ( .A(_1750_), .B(concatenador_count_0_bF_buf8), .C(_1751_), .Y(_1752_) );
	MUX2X1 MUX2X1_107 ( .A(_1752_), .B(_1749_), .S(concatenador_count_1_bF_buf0), .Y(_1753_) );
	MUX2X1 MUX2X1_108 ( .A(_1746_), .B(_1753_), .S(_1380__bF_buf5), .Y(_1754_) );
	MUX2X1 MUX2X1_109 ( .A(_1754_), .B(_1740_), .S(_1379__bF_buf0), .Y(_1755_) );
	OR2X2 OR2X2_29 ( .A(_1755_), .B(_1371_), .Y(_1756_) );
	NAND3X1 NAND3X1_83 ( .A(_1696_), .B(_1725_), .C(_1756_), .Y(_1757_) );
	INVX1 INVX1_423 ( .A(_1696_), .Y(_1758_) );
	MUX2X1 MUX2X1_110 ( .A(_1755_), .B(_1724_), .S(_1372_), .Y(_1759_) );
	NAND2X1 NAND2X1_199 ( .A(_1758_), .B(_1759_), .Y(_1760_) );
	NAND3X1 NAND3X1_84 ( .A(_1760_), .B(_1691_), .C(_1757_), .Y(_1761_) );
	AOI21X1 AOI21X1_313 ( .A(_1600_), .B(_1659_), .C(_1599_), .Y(_1762_) );
	NOR2X1 NOR2X1_144 ( .A(_1758_), .B(_1759_), .Y(_1763_) );
	AND2X2 AND2X2_44 ( .A(_1759_), .B(_1758_), .Y(_1764_) );
	OAI21X1 OAI21X1_460 ( .A(_1764_), .B(_1763_), .C(_1762_), .Y(_1765_) );
	NAND2X1 NAND2X1_200 ( .A(_1761_), .B(_1765_), .Y(_1766_) );
	OAI21X1 OAI21X1_461 ( .A(_1662_), .B(_1663_), .C(_1581_), .Y(_1767_) );
	OAI21X1 OAI21X1_462 ( .A(_1590_), .B(_1767_), .C(_1664_), .Y(_1768_) );
	AND2X2 AND2X2_45 ( .A(_1768_), .B(_1766_), .Y(_1769_) );
	OAI21X1 OAI21X1_463 ( .A(_1768_), .B(_1766_), .C(_1518_), .Y(_1770_) );
	AOI21X1 AOI21X1_314 ( .A(micro_hash_synth_c_4_), .B(_1366_), .C(_1205__bF_buf2), .Y(_1771_) );
	OAI21X1 OAI21X1_464 ( .A(_1769_), .B(_1770_), .C(_1771_), .Y(_930__4_) );
	OAI21X1 OAI21X1_465 ( .A(_1768_), .B(_1766_), .C(_1761_), .Y(_1772_) );
	AOI21X1 AOI21X1_315 ( .A(_1758_), .B(_1759_), .C(_1694_), .Y(_1773_) );
	XOR2X1 XOR2X1_30 ( .A(micro_hash_synth_k_5_), .B(micro_hash_synth_x_5_), .Y(_1774_) );
	MUX2X1 MUX2X1_111 ( .A(micro_hash_synth_W_31__5_), .B(micro_hash_synth_W_30__5_), .S(concatenador_count_0_bF_buf7), .Y(_1775_) );
	MUX2X1 MUX2X1_112 ( .A(micro_hash_synth_W_29__5_), .B(micro_hash_synth_W_28__5_), .S(concatenador_count_0_bF_buf6), .Y(_1776_) );
	MUX2X1 MUX2X1_113 ( .A(_1776_), .B(_1775_), .S(concatenador_count_1_bF_buf6), .Y(_1777_) );
	NOR2X1 NOR2X1_145 ( .A(_1373__bF_buf0), .B(_1777_), .Y(_1778_) );
	MUX2X1 MUX2X1_114 ( .A(micro_hash_synth_W_27__5_), .B(micro_hash_synth_W_26__5_), .S(concatenador_count_0_bF_buf5), .Y(_1779_) );
	MUX2X1 MUX2X1_115 ( .A(micro_hash_synth_W_25__5_), .B(micro_hash_synth_W_24__5_), .S(concatenador_count_0_bF_buf4), .Y(_1780_) );
	MUX2X1 MUX2X1_116 ( .A(_1780_), .B(_1779_), .S(concatenador_count_1_bF_buf5), .Y(_1781_) );
	OAI21X1 OAI21X1_466 ( .A(_1781_), .B(_1380__bF_buf4), .C(_1379__bF_buf3), .Y(_1782_) );
	MUX2X1 MUX2X1_117 ( .A(micro_hash_synth_W_23__5_), .B(micro_hash_synth_W_22__5_), .S(concatenador_count_0_bF_buf3), .Y(_1783_) );
	MUX2X1 MUX2X1_118 ( .A(micro_hash_synth_W_21__5_), .B(micro_hash_synth_W_20__5_), .S(concatenador_count_0_bF_buf2), .Y(_1784_) );
	MUX2X1 MUX2X1_119 ( .A(_1784_), .B(_1783_), .S(concatenador_count_1_bF_buf4), .Y(_1785_) );
	NOR2X1 NOR2X1_146 ( .A(_1373__bF_buf3), .B(_1785_), .Y(_1786_) );
	MUX2X1 MUX2X1_120 ( .A(micro_hash_synth_W_19__5_), .B(micro_hash_synth_W_18__5_), .S(concatenador_count_0_bF_buf1), .Y(_1787_) );
	MUX2X1 MUX2X1_121 ( .A(micro_hash_synth_W_17__5_), .B(micro_hash_synth_W_16__5_), .S(concatenador_count_0_bF_buf0), .Y(_1788_) );
	MUX2X1 MUX2X1_122 ( .A(_1788_), .B(_1787_), .S(concatenador_count_1_bF_buf3), .Y(_1789_) );
	OAI21X1 OAI21X1_467 ( .A(_1789_), .B(_1380__bF_buf3), .C(_1389_), .Y(_1790_) );
	OAI22X1 OAI22X1_70 ( .A(_1782_), .B(_1778_), .C(_1786_), .D(_1790_), .Y(_1791_) );
	MUX2X1 MUX2X1_123 ( .A(micro_hash_synth_W_15__5_), .B(micro_hash_synth_W_14__5_), .S(concatenador_count_0_bF_buf11), .Y(_1792_) );
	MUX2X1 MUX2X1_124 ( .A(micro_hash_synth_W_13__5_), .B(micro_hash_synth_W_12__5_), .S(concatenador_count_0_bF_buf10), .Y(_1793_) );
	MUX2X1 MUX2X1_125 ( .A(_1793_), .B(_1792_), .S(concatenador_count_1_bF_buf2), .Y(_1794_) );
	NOR2X1 NOR2X1_147 ( .A(_1373__bF_buf2), .B(_1794_), .Y(_1795_) );
	MUX2X1 MUX2X1_126 ( .A(micro_hash_synth_W_11__5_), .B(micro_hash_synth_W_10__5_), .S(concatenador_count_0_bF_buf9), .Y(_1796_) );
	MUX2X1 MUX2X1_127 ( .A(micro_hash_synth_W_9__5_), .B(micro_hash_synth_W_8__5_), .S(concatenador_count_0_bF_buf8), .Y(_1797_) );
	MUX2X1 MUX2X1_128 ( .A(_1797_), .B(_1796_), .S(concatenador_count_1_bF_buf1), .Y(_1798_) );
	OAI21X1 OAI21X1_468 ( .A(_1798_), .B(_1380__bF_buf2), .C(_1379__bF_buf2), .Y(_1799_) );
	MUX2X1 MUX2X1_129 ( .A(micro_hash_synth_W_7__5_), .B(micro_hash_synth_W_6__5_), .S(concatenador_count_0_bF_buf7), .Y(_1800_) );
	MUX2X1 MUX2X1_130 ( .A(micro_hash_synth_W_5__5_), .B(micro_hash_synth_W_4__5_), .S(concatenador_count_0_bF_buf6), .Y(_1801_) );
	MUX2X1 MUX2X1_131 ( .A(_1801_), .B(_1800_), .S(concatenador_count_1_bF_buf0), .Y(_1802_) );
	NOR2X1 NOR2X1_148 ( .A(_1373__bF_buf1), .B(_1802_), .Y(_1803_) );
	MUX2X1 MUX2X1_132 ( .A(micro_hash_synth_W_3__5_), .B(micro_hash_synth_W_2__5_), .S(concatenador_count_0_bF_buf5), .Y(_1804_) );
	MUX2X1 MUX2X1_133 ( .A(micro_hash_synth_W_1__5_), .B(micro_hash_synth_W_0__5_), .S(concatenador_count_0_bF_buf4), .Y(_1805_) );
	MUX2X1 MUX2X1_134 ( .A(_1805_), .B(_1804_), .S(concatenador_count_1_bF_buf6), .Y(_1806_) );
	OAI21X1 OAI21X1_469 ( .A(_1806_), .B(_1380__bF_buf1), .C(_1389_), .Y(_1807_) );
	OAI22X1 OAI22X1_71 ( .A(_1799_), .B(_1795_), .C(_1803_), .D(_1807_), .Y(_1808_) );
	MUX2X1 MUX2X1_135 ( .A(_1808_), .B(_1791_), .S(_1372_), .Y(_1809_) );
	XNOR2X1 XNOR2X1_26 ( .A(_1809_), .B(_1774_), .Y(_1810_) );
	XNOR2X1 XNOR2X1_27 ( .A(_1810_), .B(_1773_), .Y(_1811_) );
	XNOR2X1 XNOR2X1_28 ( .A(_1772_), .B(_1811_), .Y(_1812_) );
	AOI21X1 AOI21X1_316 ( .A(micro_hash_synth_c_5_), .B(_1366_), .C(_1205__bF_buf1), .Y(_1813_) );
	OAI21X1 OAI21X1_470 ( .A(_1812_), .B(_1522_), .C(_1813_), .Y(_930__5_) );
	NAND3X1 NAND3X1_85 ( .A(_1761_), .B(_1765_), .C(_1811_), .Y(_1814_) );
	INVX1 INVX1_424 ( .A(_1774_), .Y(_1815_) );
	NAND2X1 NAND2X1_201 ( .A(_1815_), .B(_1809_), .Y(_1816_) );
	OR2X2 OR2X2_30 ( .A(_1809_), .B(_1815_), .Y(_1817_) );
	NAND2X1 NAND2X1_202 ( .A(_1816_), .B(_1817_), .Y(_1818_) );
	NOR2X1 NOR2X1_149 ( .A(_1773_), .B(_1818_), .Y(_1819_) );
	AOI21X1 AOI21X1_317 ( .A(_1773_), .B(_1818_), .C(_1761_), .Y(_1820_) );
	NOR2X1 NOR2X1_150 ( .A(_1819_), .B(_1820_), .Y(_1821_) );
	OAI21X1 OAI21X1_471 ( .A(_1768_), .B(_1814_), .C(_1821_), .Y(_1822_) );
	INVX1 INVX1_425 ( .A(micro_hash_synth_x_5_), .Y(_1823_) );
	OAI21X1 OAI21X1_472 ( .A(_1365_), .B(_1823_), .C(_1817_), .Y(_1824_) );
	XOR2X1 XOR2X1_31 ( .A(micro_hash_synth_k_6_), .B(micro_hash_synth_x_6_), .Y(_1825_) );
	AOI22X1 AOI22X1_30 ( .A(micro_hash_synth_W_18__6_), .B(_2470__bF_buf3), .C(_1549__bF_buf2), .D(micro_hash_synth_W_19__6_), .Y(_1826_) );
	AOI22X1 AOI22X1_31 ( .A(micro_hash_synth_W_17__6_), .B(_1547__bF_buf2), .C(_2609__bF_buf1), .D(micro_hash_synth_W_16__6_), .Y(_1827_) );
	AOI21X1 AOI21X1_318 ( .A(_1826_), .B(_1827_), .C(_1380__bF_buf0), .Y(_1828_) );
	AOI22X1 AOI22X1_32 ( .A(micro_hash_synth_W_22__6_), .B(_2470__bF_buf2), .C(_1549__bF_buf1), .D(micro_hash_synth_W_23__6_), .Y(_1829_) );
	AOI22X1 AOI22X1_33 ( .A(micro_hash_synth_W_21__6_), .B(_1547__bF_buf1), .C(_2609__bF_buf0), .D(micro_hash_synth_W_20__6_), .Y(_1830_) );
	NAND2X1 NAND2X1_203 ( .A(_1829_), .B(_1830_), .Y(_1831_) );
	AOI21X1 AOI21X1_319 ( .A(_1380__bF_buf6), .B(_1831_), .C(_1828_), .Y(_1832_) );
	AOI22X1 AOI22X1_34 ( .A(micro_hash_synth_W_30__6_), .B(_2470__bF_buf1), .C(_1549__bF_buf0), .D(micro_hash_synth_W_31__6_), .Y(_1833_) );
	AOI22X1 AOI22X1_35 ( .A(micro_hash_synth_W_29__6_), .B(_1547__bF_buf0), .C(_2609__bF_buf3), .D(micro_hash_synth_W_28__6_), .Y(_1834_) );
	NAND2X1 NAND2X1_204 ( .A(_1833_), .B(_1834_), .Y(_1835_) );
	NOR2X1 NOR2X1_151 ( .A(_1373__bF_buf0), .B(_1835_), .Y(_1836_) );
	AOI22X1 AOI22X1_36 ( .A(micro_hash_synth_W_26__6_), .B(_2470__bF_buf0), .C(_1549__bF_buf3), .D(micro_hash_synth_W_27__6_), .Y(_1837_) );
	AOI22X1 AOI22X1_37 ( .A(micro_hash_synth_W_25__6_), .B(_1547__bF_buf3), .C(_2609__bF_buf2), .D(micro_hash_synth_W_24__6_), .Y(_1838_) );
	NAND2X1 NAND2X1_205 ( .A(_1837_), .B(_1838_), .Y(_1839_) );
	OAI21X1 OAI21X1_473 ( .A(_1839_), .B(_1380__bF_buf5), .C(_1379__bF_buf1), .Y(_1840_) );
	OAI22X1 OAI22X1_72 ( .A(_1840_), .B(_1836_), .C(_1832_), .D(_1379__bF_buf0), .Y(_1841_) );
	AOI22X1 AOI22X1_38 ( .A(micro_hash_synth_W_6__6_), .B(_2470__bF_buf3), .C(_1549__bF_buf2), .D(micro_hash_synth_W_7__6_), .Y(_1842_) );
	AOI22X1 AOI22X1_39 ( .A(micro_hash_synth_W_5__6_), .B(_1547__bF_buf2), .C(_2609__bF_buf1), .D(micro_hash_synth_W_4__6_), .Y(_1843_) );
	AOI21X1 AOI21X1_320 ( .A(_1842_), .B(_1843_), .C(_1373__bF_buf3), .Y(_1844_) );
	AOI22X1 AOI22X1_40 ( .A(micro_hash_synth_W_2__6_), .B(_2470__bF_buf2), .C(_1549__bF_buf1), .D(micro_hash_synth_W_3__6_), .Y(_1845_) );
	AOI22X1 AOI22X1_41 ( .A(micro_hash_synth_W_1__6_), .B(_1547__bF_buf1), .C(_2609__bF_buf0), .D(micro_hash_synth_W_0__6_), .Y(_1846_) );
	NAND2X1 NAND2X1_206 ( .A(_1845_), .B(_1846_), .Y(_1847_) );
	AOI21X1 AOI21X1_321 ( .A(_1373__bF_buf2), .B(_1847_), .C(_1844_), .Y(_1848_) );
	AOI22X1 AOI22X1_42 ( .A(micro_hash_synth_W_14__6_), .B(_2470__bF_buf1), .C(_1549__bF_buf0), .D(micro_hash_synth_W_15__6_), .Y(_1849_) );
	AOI22X1 AOI22X1_43 ( .A(micro_hash_synth_W_13__6_), .B(_1547__bF_buf0), .C(_2609__bF_buf3), .D(micro_hash_synth_W_12__6_), .Y(_1850_) );
	NAND2X1 NAND2X1_207 ( .A(_1849_), .B(_1850_), .Y(_1851_) );
	NOR2X1 NOR2X1_152 ( .A(_1373__bF_buf1), .B(_1851_), .Y(_1852_) );
	AOI22X1 AOI22X1_44 ( .A(micro_hash_synth_W_10__6_), .B(_2470__bF_buf0), .C(_1549__bF_buf3), .D(micro_hash_synth_W_11__6_), .Y(_1853_) );
	AOI22X1 AOI22X1_45 ( .A(micro_hash_synth_W_9__6_), .B(_1547__bF_buf3), .C(_2609__bF_buf2), .D(micro_hash_synth_W_8__6_), .Y(_1854_) );
	NAND2X1 NAND2X1_208 ( .A(_1853_), .B(_1854_), .Y(_1855_) );
	OAI21X1 OAI21X1_474 ( .A(_1855_), .B(_1380__bF_buf4), .C(_1379__bF_buf3), .Y(_1856_) );
	OAI22X1 OAI22X1_73 ( .A(_1856_), .B(_1852_), .C(_1848_), .D(_1379__bF_buf2), .Y(_1857_) );
	MUX2X1 MUX2X1_136 ( .A(_1857_), .B(_1841_), .S(_1372_), .Y(_1858_) );
	XNOR2X1 XNOR2X1_29 ( .A(_1858_), .B(_1825_), .Y(_1859_) );
	AND2X2 AND2X2_46 ( .A(_1859_), .B(_1824_), .Y(_1860_) );
	NOR2X1 NOR2X1_153 ( .A(_1824_), .B(_1859_), .Y(_1861_) );
	NOR2X1 NOR2X1_154 ( .A(_1861_), .B(_1860_), .Y(_1862_) );
	NOR2X1 NOR2X1_155 ( .A(_1862_), .B(_1822_), .Y(_1863_) );
	NOR2X1 NOR2X1_156 ( .A(_1584_), .B(_1583_), .Y(_1864_) );
	AOI22X1 AOI22X1_46 ( .A(_1596_), .B(_1660_), .C(_1864_), .D(_1524_), .Y(_1865_) );
	OAI21X1 OAI21X1_475 ( .A(_1586_), .B(_1519_), .C(_1865_), .Y(_1866_) );
	OAI21X1 OAI21X1_476 ( .A(_1694_), .B(_1764_), .C(_1818_), .Y(_1867_) );
	NAND2X1 NAND2X1_209 ( .A(_1773_), .B(_1810_), .Y(_1868_) );
	AOI21X1 AOI21X1_322 ( .A(_1867_), .B(_1868_), .C(_1766_), .Y(_1869_) );
	NAND3X1 NAND3X1_86 ( .A(_1664_), .B(_1866_), .C(_1869_), .Y(_1870_) );
	INVX1 INVX1_426 ( .A(_1862_), .Y(_1871_) );
	AOI21X1 AOI21X1_323 ( .A(_1821_), .B(_1870_), .C(_1871_), .Y(_1872_) );
	OR2X2 OR2X2_31 ( .A(_1872_), .B(_1522_), .Y(_1873_) );
	AOI21X1 AOI21X1_324 ( .A(micro_hash_synth_c_6_), .B(_1366_), .C(_1205__bF_buf0), .Y(_1874_) );
	OAI21X1 OAI21X1_477 ( .A(_1873_), .B(_1863_), .C(_1874_), .Y(_930__6_) );
	NAND2X1 NAND2X1_210 ( .A(micro_hash_synth_k_6_), .B(micro_hash_synth_x_6_), .Y(_1875_) );
	INVX1 INVX1_427 ( .A(_1825_), .Y(_1876_) );
	OAI21X1 OAI21X1_478 ( .A(_1858_), .B(_1876_), .C(_1875_), .Y(_1877_) );
	XOR2X1 XOR2X1_32 ( .A(micro_hash_synth_k_7_), .B(micro_hash_synth_x_7_), .Y(_1878_) );
	AOI22X1 AOI22X1_47 ( .A(micro_hash_synth_W_26__7_), .B(_2470__bF_buf3), .C(_1549__bF_buf2), .D(micro_hash_synth_W_27__7_), .Y(_1879_) );
	AOI22X1 AOI22X1_48 ( .A(micro_hash_synth_W_25__7_), .B(_1547__bF_buf2), .C(_2609__bF_buf1), .D(micro_hash_synth_W_24__7_), .Y(_1880_) );
	AOI21X1 AOI21X1_325 ( .A(_1879_), .B(_1880_), .C(_1380__bF_buf3), .Y(_1881_) );
	AOI22X1 AOI22X1_49 ( .A(micro_hash_synth_W_30__7_), .B(_2470__bF_buf2), .C(_1549__bF_buf1), .D(micro_hash_synth_W_31__7_), .Y(_1882_) );
	AOI22X1 AOI22X1_50 ( .A(micro_hash_synth_W_29__7_), .B(_1547__bF_buf1), .C(_2609__bF_buf0), .D(micro_hash_synth_W_28__7_), .Y(_1883_) );
	NAND2X1 NAND2X1_211 ( .A(_1882_), .B(_1883_), .Y(_1884_) );
	AOI21X1 AOI21X1_326 ( .A(_1380__bF_buf2), .B(_1884_), .C(_1881_), .Y(_1885_) );
	AOI22X1 AOI22X1_51 ( .A(micro_hash_synth_W_22__7_), .B(_2470__bF_buf1), .C(_1549__bF_buf0), .D(micro_hash_synth_W_23__7_), .Y(_1886_) );
	AOI22X1 AOI22X1_52 ( .A(micro_hash_synth_W_21__7_), .B(_1547__bF_buf0), .C(_2609__bF_buf3), .D(micro_hash_synth_W_20__7_), .Y(_1887_) );
	NAND2X1 NAND2X1_212 ( .A(_1886_), .B(_1887_), .Y(_1888_) );
	NOR2X1 NOR2X1_157 ( .A(_1373__bF_buf0), .B(_1888_), .Y(_1889_) );
	AOI22X1 AOI22X1_53 ( .A(micro_hash_synth_W_17__7_), .B(_1547__bF_buf3), .C(_2609__bF_buf2), .D(micro_hash_synth_W_16__7_), .Y(_1890_) );
	AOI22X1 AOI22X1_54 ( .A(micro_hash_synth_W_18__7_), .B(_2470__bF_buf0), .C(_1549__bF_buf3), .D(micro_hash_synth_W_19__7_), .Y(_1891_) );
	NAND2X1 NAND2X1_213 ( .A(_1891_), .B(_1890_), .Y(_1892_) );
	OAI21X1 OAI21X1_479 ( .A(_1892_), .B(_1380__bF_buf1), .C(_1389_), .Y(_1893_) );
	OAI22X1 OAI22X1_74 ( .A(_1893_), .B(_1889_), .C(_1885_), .D(_1389_), .Y(_1894_) );
	AOI22X1 AOI22X1_55 ( .A(micro_hash_synth_W_14__7_), .B(_2470__bF_buf3), .C(_1549__bF_buf2), .D(micro_hash_synth_W_15__7_), .Y(_1895_) );
	AOI22X1 AOI22X1_56 ( .A(micro_hash_synth_W_13__7_), .B(_1547__bF_buf2), .C(_2609__bF_buf1), .D(micro_hash_synth_W_12__7_), .Y(_1896_) );
	AOI21X1 AOI21X1_327 ( .A(_1895_), .B(_1896_), .C(_1373__bF_buf3), .Y(_1897_) );
	AOI22X1 AOI22X1_57 ( .A(micro_hash_synth_W_10__7_), .B(_2470__bF_buf2), .C(_1549__bF_buf1), .D(micro_hash_synth_W_11__7_), .Y(_1898_) );
	AOI22X1 AOI22X1_58 ( .A(micro_hash_synth_W_9__7_), .B(_1547__bF_buf1), .C(_2609__bF_buf0), .D(micro_hash_synth_W_8__7_), .Y(_1899_) );
	NAND2X1 NAND2X1_214 ( .A(_1898_), .B(_1899_), .Y(_1900_) );
	AOI21X1 AOI21X1_328 ( .A(_1373__bF_buf2), .B(_1900_), .C(_1897_), .Y(_1901_) );
	AOI22X1 AOI22X1_59 ( .A(micro_hash_synth_W_6__7_), .B(_2470__bF_buf1), .C(_1549__bF_buf0), .D(micro_hash_synth_W_7__7_), .Y(_1902_) );
	AOI22X1 AOI22X1_60 ( .A(micro_hash_synth_W_5__7_), .B(_1547__bF_buf0), .C(_2609__bF_buf3), .D(micro_hash_synth_W_4__7_), .Y(_1903_) );
	NAND2X1 NAND2X1_215 ( .A(_1902_), .B(_1903_), .Y(_1904_) );
	NOR2X1 NOR2X1_158 ( .A(_1373__bF_buf1), .B(_1904_), .Y(_1905_) );
	AOI22X1 AOI22X1_61 ( .A(micro_hash_synth_W_1__7_), .B(_1547__bF_buf3), .C(_2609__bF_buf2), .D(micro_hash_synth_W_0__7_), .Y(_1906_) );
	AOI22X1 AOI22X1_62 ( .A(micro_hash_synth_W_2__7_), .B(_2470__bF_buf0), .C(_1549__bF_buf3), .D(micro_hash_synth_W_3__7_), .Y(_1907_) );
	NAND2X1 NAND2X1_216 ( .A(_1907_), .B(_1906_), .Y(_1908_) );
	OAI21X1 OAI21X1_480 ( .A(_1908_), .B(_1380__bF_buf0), .C(_1389_), .Y(_1909_) );
	OAI22X1 OAI22X1_75 ( .A(_1909_), .B(_1905_), .C(_1901_), .D(_1389_), .Y(_1910_) );
	MUX2X1 MUX2X1_137 ( .A(_1910_), .B(_1894_), .S(_1372_), .Y(_1911_) );
	XOR2X1 XOR2X1_33 ( .A(_1911_), .B(_1878_), .Y(_1912_) );
	XNOR2X1 XNOR2X1_30 ( .A(_1912_), .B(_1877_), .Y(_1913_) );
	NOR3X1 NOR3X1_3 ( .A(_1860_), .B(_1913_), .C(_1872_), .Y(_1914_) );
	AOI21X1 AOI21X1_329 ( .A(_1862_), .B(_1822_), .C(_1860_), .Y(_1915_) );
	INVX1 INVX1_428 ( .A(_1913_), .Y(_1916_) );
	OAI21X1 OAI21X1_481 ( .A(_1915_), .B(_1916_), .C(_1518_), .Y(_1917_) );
	AOI21X1 AOI21X1_330 ( .A(micro_hash_synth_c_7_), .B(_1366_), .C(_1205__bF_buf3), .Y(_1918_) );
	OAI21X1 OAI21X1_482 ( .A(_1917_), .B(_1914_), .C(_1918_), .Y(_930__7_) );
	OAI21X1 OAI21X1_483 ( .A(_1256_), .B(_1354__bF_buf3), .C(_1269__bF_buf0), .Y(_929__0_) );
	NOR2X1 NOR2X1_159 ( .A(_1262_), .B(_1356_), .Y(_929__1_) );
	AND2X2 AND2X2_47 ( .A(_1355_), .B(micro_hash_synth_b_2_), .Y(_929__2_) );
	INVX1 INVX1_429 ( .A(micro_hash_synth_b_3_), .Y(_1919_) );
	OAI21X1 OAI21X1_484 ( .A(_1919_), .B(_1354__bF_buf2), .C(_1269__bF_buf3), .Y(_929__3_) );
	OAI21X1 OAI21X1_485 ( .A(micro_hash_synth_b_4_), .B(_1354__bF_buf1), .C(_1269__bF_buf2), .Y(_1920_) );
	AOI21X1 AOI21X1_331 ( .A(_1367_), .B(_1518_), .C(_1920_), .Y(_929__4_) );
	OAI21X1 OAI21X1_486 ( .A(micro_hash_synth_b_5_), .B(_1354__bF_buf0), .C(_1269__bF_buf1), .Y(_1921_) );
	AOI21X1 AOI21X1_332 ( .A(_1208_), .B(_1518_), .C(_1921_), .Y(_929__5_) );
	OAI21X1 OAI21X1_487 ( .A(micro_hash_synth_b_6_), .B(_1354__bF_buf3), .C(_1269__bF_buf0), .Y(_1922_) );
	AOI21X1 AOI21X1_333 ( .A(_1216_), .B(_1518_), .C(_1922_), .Y(_929__6_) );
	INVX1 INVX1_430 ( .A(micro_hash_synth_c_3_), .Y(_1923_) );
	INVX1 INVX1_431 ( .A(micro_hash_synth_b_7_), .Y(_1924_) );
	AOI22X1 AOI22X1_63 ( .A(_1924_), .B(_1355_), .C(_1415_), .D(_1923_), .Y(_929__7_) );
	XNOR2X1 XNOR2X1_31 ( .A(micro_hash_synth_c_0_), .B(micro_hash_synth_b_0_), .Y(_1925_) );
	AOI21X1 AOI21X1_334 ( .A(micro_hash_synth_a_0_), .B(_1366_), .C(_1205__bF_buf2), .Y(_1926_) );
	OAI21X1 OAI21X1_488 ( .A(_1522_), .B(_1925_), .C(_1926_), .Y(_928__0_) );
	INVX2 INVX2_4 ( .A(_1415_), .Y(_1927_) );
	XNOR2X1 XNOR2X1_32 ( .A(micro_hash_synth_c_1_), .B(micro_hash_synth_b_1_), .Y(_1928_) );
	OAI22X1 OAI22X1_76 ( .A(_1310_), .B(_1356_), .C(_1927_), .D(_1928_), .Y(_928__1_) );
	NAND2X1 NAND2X1_217 ( .A(micro_hash_synth_a_2_), .B(_1355_), .Y(_1929_) );
	XNOR2X1 XNOR2X1_33 ( .A(micro_hash_synth_c_2_), .B(micro_hash_synth_b_2_), .Y(_1930_) );
	OAI21X1 OAI21X1_489 ( .A(_1927_), .B(_1930_), .C(_1929_), .Y(_928__2_) );
	INVX1 INVX1_432 ( .A(micro_hash_synth_a_3_), .Y(_1931_) );
	XNOR2X1 XNOR2X1_34 ( .A(micro_hash_synth_c_3_), .B(micro_hash_synth_b_3_), .Y(_1932_) );
	OAI22X1 OAI22X1_77 ( .A(_1931_), .B(_1356_), .C(_1927_), .D(_1932_), .Y(_928__3_) );
	NAND2X1 NAND2X1_218 ( .A(micro_hash_synth_a_4_), .B(_1355_), .Y(_1933_) );
	XNOR2X1 XNOR2X1_35 ( .A(micro_hash_synth_c_4_), .B(micro_hash_synth_b_4_), .Y(_1934_) );
	OAI21X1 OAI21X1_490 ( .A(_1927_), .B(_1934_), .C(_1933_), .Y(_928__4_) );
	NAND2X1 NAND2X1_219 ( .A(micro_hash_synth_a_5_), .B(_1355_), .Y(_1935_) );
	XNOR2X1 XNOR2X1_36 ( .A(micro_hash_synth_c_5_), .B(micro_hash_synth_b_5_), .Y(_1936_) );
	OAI21X1 OAI21X1_491 ( .A(_1927_), .B(_1936_), .C(_1935_), .Y(_928__5_) );
	XNOR2X1 XNOR2X1_37 ( .A(micro_hash_synth_c_6_), .B(micro_hash_synth_b_6_), .Y(_1937_) );
	OAI22X1 OAI22X1_78 ( .A(_1349_), .B(_1356_), .C(_1927_), .D(_1937_), .Y(_928__6_) );
	NAND2X1 NAND2X1_220 ( .A(micro_hash_synth_a_7_), .B(_1355_), .Y(_1938_) );
	XNOR2X1 XNOR2X1_38 ( .A(micro_hash_synth_c_7_), .B(micro_hash_synth_b_7_), .Y(_1939_) );
	OAI21X1 OAI21X1_492 ( .A(_1927_), .B(_1939_), .C(_1938_), .Y(_928__7_) );
	INVX1 INVX1_433 ( .A(bloque_in_0_), .Y(_1940_) );
	NOR2X1 NOR2X1_160 ( .A(_1202__bF_buf2), .B(_1940_), .Y(_933__0_) );
	INVX1 INVX1_434 ( .A(bloque_in_1_), .Y(_1941_) );
	NOR2X1 NOR2X1_161 ( .A(_1202__bF_buf1), .B(_1941_), .Y(_933__1_) );
	INVX1 INVX1_435 ( .A(bloque_in_2_), .Y(_1942_) );
	NOR2X1 NOR2X1_162 ( .A(_1202__bF_buf0), .B(_1942_), .Y(_933__2_) );
	INVX1 INVX1_436 ( .A(bloque_in_3_), .Y(_1943_) );
	NOR2X1 NOR2X1_163 ( .A(_1202__bF_buf5), .B(_1943_), .Y(_933__3_) );
	INVX1 INVX1_437 ( .A(bloque_in_4_), .Y(_1944_) );
	NOR2X1 NOR2X1_164 ( .A(_1202__bF_buf4), .B(_1944_), .Y(_933__4_) );
	INVX1 INVX1_438 ( .A(bloque_in_5_), .Y(_1945_) );
	NOR2X1 NOR2X1_165 ( .A(_1202__bF_buf3), .B(_1945_), .Y(_933__5_) );
	INVX1 INVX1_439 ( .A(bloque_in_6_), .Y(_1946_) );
	NOR2X1 NOR2X1_166 ( .A(_1202__bF_buf2), .B(_1946_), .Y(_933__6_) );
	INVX1 INVX1_440 ( .A(bloque_in_7_), .Y(_1947_) );
	NOR2X1 NOR2X1_167 ( .A(_1202__bF_buf1), .B(_1947_), .Y(_933__7_) );
	INVX1 INVX1_441 ( .A(bloque_in_8_), .Y(_1948_) );
	NOR2X1 NOR2X1_168 ( .A(_1202__bF_buf0), .B(_1948_), .Y(_933__8_) );
	INVX1 INVX1_442 ( .A(bloque_in_9_), .Y(_1949_) );
	NOR2X1 NOR2X1_169 ( .A(_1202__bF_buf5), .B(_1949_), .Y(_933__9_) );
	INVX1 INVX1_443 ( .A(bloque_in_10_), .Y(_1950_) );
	NOR2X1 NOR2X1_170 ( .A(_1202__bF_buf4), .B(_1950_), .Y(_933__10_) );
	INVX1 INVX1_444 ( .A(bloque_in_11_), .Y(_1951_) );
	NOR2X1 NOR2X1_171 ( .A(_1202__bF_buf3), .B(_1951_), .Y(_933__11_) );
	INVX1 INVX1_445 ( .A(bloque_in_12_), .Y(_1952_) );
	NOR2X1 NOR2X1_172 ( .A(_1202__bF_buf2), .B(_1952_), .Y(_933__12_) );
	INVX1 INVX1_446 ( .A(bloque_in_13_), .Y(_1953_) );
	NOR2X1 NOR2X1_173 ( .A(_1202__bF_buf1), .B(_1953_), .Y(_933__13_) );
	INVX1 INVX1_447 ( .A(bloque_in_14_), .Y(_1954_) );
	NOR2X1 NOR2X1_174 ( .A(_1202__bF_buf0), .B(_1954_), .Y(_933__14_) );
	INVX1 INVX1_448 ( .A(bloque_in_15_), .Y(_1955_) );
	NOR2X1 NOR2X1_175 ( .A(_1202__bF_buf5), .B(_1955_), .Y(_933__15_) );
	INVX1 INVX1_449 ( .A(bloque_in_16_), .Y(_1956_) );
	NOR2X1 NOR2X1_176 ( .A(_1202__bF_buf4), .B(_1956_), .Y(_933__16_) );
	INVX1 INVX1_450 ( .A(bloque_in_17_), .Y(_1957_) );
	NOR2X1 NOR2X1_177 ( .A(_1202__bF_buf3), .B(_1957_), .Y(_933__17_) );
	INVX1 INVX1_451 ( .A(bloque_in_18_), .Y(_1958_) );
	NOR2X1 NOR2X1_178 ( .A(_1202__bF_buf2), .B(_1958_), .Y(_933__18_) );
	INVX1 INVX1_452 ( .A(bloque_in_19_), .Y(_1959_) );
	NOR2X1 NOR2X1_179 ( .A(_1202__bF_buf1), .B(_1959_), .Y(_933__19_) );
	INVX1 INVX1_453 ( .A(bloque_in_20_), .Y(_1960_) );
	NOR2X1 NOR2X1_180 ( .A(_1202__bF_buf0), .B(_1960_), .Y(_933__20_) );
	INVX1 INVX1_454 ( .A(bloque_in_21_), .Y(_1961_) );
	NOR2X1 NOR2X1_181 ( .A(_1202__bF_buf5), .B(_1961_), .Y(_933__21_) );
	INVX1 INVX1_455 ( .A(bloque_in_22_), .Y(_1962_) );
	NOR2X1 NOR2X1_182 ( .A(_1202__bF_buf4), .B(_1962_), .Y(_933__22_) );
	INVX1 INVX1_456 ( .A(bloque_in_23_), .Y(_1963_) );
	NOR2X1 NOR2X1_183 ( .A(_1202__bF_buf3), .B(_1963_), .Y(_933__23_) );
	INVX1 INVX1_457 ( .A(bloque_in_24_), .Y(_1964_) );
	NOR2X1 NOR2X1_184 ( .A(_1202__bF_buf2), .B(_1964_), .Y(_933__24_) );
	INVX1 INVX1_458 ( .A(bloque_in_25_), .Y(_1965_) );
	NOR2X1 NOR2X1_185 ( .A(_1202__bF_buf1), .B(_1965_), .Y(_933__25_) );
	INVX1 INVX1_459 ( .A(bloque_in_26_), .Y(_1966_) );
	NOR2X1 NOR2X1_186 ( .A(_1202__bF_buf0), .B(_1966_), .Y(_933__26_) );
	INVX1 INVX1_460 ( .A(bloque_in_27_), .Y(_1967_) );
	NOR2X1 NOR2X1_187 ( .A(_1202__bF_buf5), .B(_1967_), .Y(_933__27_) );
	INVX1 INVX1_461 ( .A(bloque_in_28_), .Y(_1968_) );
	NOR2X1 NOR2X1_188 ( .A(_1202__bF_buf4), .B(_1968_), .Y(_933__28_) );
	INVX1 INVX1_462 ( .A(bloque_in_29_), .Y(_1969_) );
	NOR2X1 NOR2X1_189 ( .A(_1202__bF_buf3), .B(_1969_), .Y(_933__29_) );
	INVX1 INVX1_463 ( .A(bloque_in_30_), .Y(_1970_) );
	NOR2X1 NOR2X1_190 ( .A(_1202__bF_buf2), .B(_1970_), .Y(_933__30_) );
	INVX1 INVX1_464 ( .A(bloque_in_31_), .Y(_1971_) );
	NOR2X1 NOR2X1_191 ( .A(_1202__bF_buf1), .B(_1971_), .Y(_933__31_) );
	NAND2X1 NAND2X1_221 ( .A(_2462_), .B(_1354__bF_buf2), .Y(_1972_) );
	NAND2X1 NAND2X1_222 ( .A(concatenador_count_0_bF_buf3), .B(_1366_), .Y(_1973_) );
	AOI21X1 AOI21X1_335 ( .A(_1972_), .B(_1973_), .C(_1254_), .Y(_931__0_) );
	OAI21X1 OAI21X1_493 ( .A(_2609__bF_buf1), .B(_1549__bF_buf2), .C(_1518_), .Y(_1974_) );
	AOI21X1 AOI21X1_336 ( .A(concatenador_count_1_bF_buf5), .B(_1366_), .C(_2472_), .Y(_1975_) );
	AOI21X1 AOI21X1_337 ( .A(_1974_), .B(_1975_), .C(_1254_), .Y(_931__1_) );
	INVX1 INVX1_465 ( .A(concatenador_count_2_), .Y(_1976_) );
	NAND2X1 NAND2X1_223 ( .A(_2610_), .B(_1547__bF_buf2), .Y(_1977_) );
	XNOR2X1 XNOR2X1_39 ( .A(_1977_), .B(_1976_), .Y(_1978_) );
	NOR2X1 NOR2X1_192 ( .A(_1978_), .B(_1254_), .Y(_931__2_) );
	NAND2X1 NAND2X1_224 ( .A(concatenador_count_3_), .B(concatenador_count_2_), .Y(_1979_) );
	NOR2X1 NOR2X1_193 ( .A(_1433_), .B(_1979_), .Y(_1980_) );
	NAND2X1 NAND2X1_225 ( .A(_1980_), .B(_1518_), .Y(_1981_) );
	INVX1 INVX1_466 ( .A(concatenador_count_3_), .Y(_1982_) );
	OAI21X1 OAI21X1_494 ( .A(_1977_), .B(_1976_), .C(_1982_), .Y(_1983_) );
	NAND2X1 NAND2X1_226 ( .A(_1983_), .B(_1981_), .Y(_1984_) );
	NOR2X1 NOR2X1_194 ( .A(_1254_), .B(_1984_), .Y(_931__3_) );
	NAND2X1 NAND2X1_227 ( .A(concatenador_count_4_), .B(_1980_), .Y(_1985_) );
	OAI21X1 OAI21X1_495 ( .A(concatenador_count_5_), .B(_1985_), .C(_1253_), .Y(_1986_) );
	AOI21X1 AOI21X1_338 ( .A(_1360_), .B(_1981_), .C(_1986_), .Y(_931__4_) );
	AOI21X1 AOI21X1_339 ( .A(_2610_), .B(_1985_), .C(_1254_), .Y(_931__5_) );
	NOR2X1 NOR2X1_195 ( .A(micro_hash_synth_x_0_), .B(_1354__bF_buf1), .Y(_1987_) );
	NAND2X1 NAND2X1_228 ( .A(_1256_), .B(_1306_), .Y(_1988_) );
	OAI21X1 OAI21X1_496 ( .A(_1366_), .B(_1988_), .C(_1363_), .Y(_1989_) );
	NOR2X1 NOR2X1_196 ( .A(concatenador_count_5_), .B(_1361_), .Y(_1990_) );
	XOR2X1 XOR2X1_34 ( .A(micro_hash_synth_b_0_), .B(micro_hash_synth_a_0_), .Y(_1991_) );
	NAND3X1 NAND3X1_87 ( .A(_1990_), .B(_1991_), .C(_1269__bF_buf3), .Y(_1992_) );
	OAI21X1 OAI21X1_497 ( .A(_1989_), .B(_1987_), .C(_1992_), .Y(_934__0_) );
	OAI21X1 OAI21X1_498 ( .A(micro_hash_synth_b_1_), .B(micro_hash_synth_a_1_), .C(_1354__bF_buf0), .Y(_1993_) );
	OAI21X1 OAI21X1_499 ( .A(_1419_), .B(_1354__bF_buf3), .C(_1993_), .Y(_1994_) );
	OAI21X1 OAI21X1_500 ( .A(concatenador_count_5_), .B(_1361_), .C(_1994_), .Y(_1995_) );
	XOR2X1 XOR2X1_35 ( .A(micro_hash_synth_b_1_), .B(micro_hash_synth_a_1_), .Y(_1996_) );
	NAND3X1 NAND3X1_88 ( .A(_1990_), .B(_1996_), .C(_1269__bF_buf2), .Y(_1997_) );
	OAI21X1 OAI21X1_501 ( .A(_1995_), .B(_1202__bF_buf0), .C(_1997_), .Y(_934__1_) );
	OAI21X1 OAI21X1_502 ( .A(micro_hash_synth_b_2_), .B(micro_hash_synth_a_2_), .C(_1354__bF_buf2), .Y(_1998_) );
	OAI21X1 OAI21X1_503 ( .A(_1595_), .B(_1354__bF_buf1), .C(_1998_), .Y(_1999_) );
	OAI21X1 OAI21X1_504 ( .A(concatenador_count_5_), .B(_1361_), .C(_1999_), .Y(_2000_) );
	XOR2X1 XOR2X1_36 ( .A(micro_hash_synth_b_2_), .B(micro_hash_synth_a_2_), .Y(_2001_) );
	NAND3X1 NAND3X1_89 ( .A(_1990_), .B(_2001_), .C(_1269__bF_buf1), .Y(_2002_) );
	OAI21X1 OAI21X1_505 ( .A(_2000_), .B(_1202__bF_buf5), .C(_2002_), .Y(_934__2_) );
	NOR2X1 NOR2X1_197 ( .A(micro_hash_synth_b_3_), .B(micro_hash_synth_a_3_), .Y(_2003_) );
	NOR2X1 NOR2X1_198 ( .A(_2003_), .B(_1366_), .Y(_2004_) );
	AOI21X1 AOI21X1_340 ( .A(micro_hash_synth_x_3_), .B(_1366_), .C(_2004_), .Y(_2005_) );
	NOR2X1 NOR2X1_199 ( .A(_1919_), .B(_1931_), .Y(_2006_) );
	OAI21X1 OAI21X1_506 ( .A(_2003_), .B(_2006_), .C(_1269__bF_buf0), .Y(_2007_) );
	OAI21X1 OAI21X1_507 ( .A(_1202__bF_buf4), .B(_1990_), .C(_2007_), .Y(_2008_) );
	OAI21X1 OAI21X1_508 ( .A(_2005_), .B(_1990_), .C(_2008_), .Y(_934__3_) );
	OAI21X1 OAI21X1_509 ( .A(micro_hash_synth_b_4_), .B(micro_hash_synth_a_4_), .C(_1354__bF_buf0), .Y(_2009_) );
	OAI21X1 OAI21X1_510 ( .A(_1692_), .B(_1354__bF_buf3), .C(_2009_), .Y(_2010_) );
	OAI21X1 OAI21X1_511 ( .A(concatenador_count_5_), .B(_1361_), .C(_2010_), .Y(_2011_) );
	XOR2X1 XOR2X1_37 ( .A(micro_hash_synth_b_4_), .B(micro_hash_synth_a_4_), .Y(_2012_) );
	NAND3X1 NAND3X1_90 ( .A(_1990_), .B(_2012_), .C(_1269__bF_buf3), .Y(_2013_) );
	OAI21X1 OAI21X1_512 ( .A(_2011_), .B(_1202__bF_buf3), .C(_2013_), .Y(_934__4_) );
	OAI21X1 OAI21X1_513 ( .A(micro_hash_synth_b_5_), .B(micro_hash_synth_a_5_), .C(_1354__bF_buf2), .Y(_2014_) );
	OAI21X1 OAI21X1_514 ( .A(_1823_), .B(_1354__bF_buf1), .C(_2014_), .Y(_2015_) );
	OAI21X1 OAI21X1_515 ( .A(concatenador_count_5_), .B(_1361_), .C(_2015_), .Y(_2016_) );
	XOR2X1 XOR2X1_38 ( .A(micro_hash_synth_b_5_), .B(micro_hash_synth_a_5_), .Y(_2017_) );
	NAND3X1 NAND3X1_91 ( .A(_1990_), .B(_2017_), .C(_1269__bF_buf2), .Y(_2018_) );
	OAI21X1 OAI21X1_516 ( .A(_2016_), .B(_1202__bF_buf2), .C(_2018_), .Y(_934__5_) );
	NOR2X1 NOR2X1_200 ( .A(micro_hash_synth_b_6_), .B(micro_hash_synth_a_6_), .Y(_2019_) );
	AOI21X1 AOI21X1_341 ( .A(_2019_), .B(_1354__bF_buf0), .C(_1990_), .Y(_2020_) );
	OAI21X1 OAI21X1_517 ( .A(micro_hash_synth_x_6_), .B(_1354__bF_buf3), .C(_2020_), .Y(_2021_) );
	XOR2X1 XOR2X1_39 ( .A(micro_hash_synth_b_6_), .B(micro_hash_synth_a_6_), .Y(_2022_) );
	NAND3X1 NAND3X1_92 ( .A(_1990_), .B(_2022_), .C(_1269__bF_buf1), .Y(_2023_) );
	OAI21X1 OAI21X1_518 ( .A(_2021_), .B(_1202__bF_buf1), .C(_2023_), .Y(_934__6_) );
	NOR2X1 NOR2X1_201 ( .A(micro_hash_synth_b_7_), .B(micro_hash_synth_a_7_), .Y(_2024_) );
	NAND2X1 NAND2X1_229 ( .A(_2024_), .B(_1354__bF_buf2), .Y(_2025_) );
	OAI21X1 OAI21X1_519 ( .A(micro_hash_synth_x_7_), .B(_1354__bF_buf1), .C(_2025_), .Y(_2026_) );
	AND2X2 AND2X2_48 ( .A(micro_hash_synth_b_7_), .B(micro_hash_synth_a_7_), .Y(_2027_) );
	OAI21X1 OAI21X1_520 ( .A(_2024_), .B(_2027_), .C(_1269__bF_buf0), .Y(_2028_) );
	OAI21X1 OAI21X1_521 ( .A(_1202__bF_buf0), .B(_1990_), .C(_2028_), .Y(_2029_) );
	OAI21X1 OAI21X1_522 ( .A(_2026_), .B(_1990_), .C(_2029_), .Y(_934__7_) );
	INVX1 INVX1_467 ( .A(micro_hash_synth_W_3__0_), .Y(_2030_) );
	OAI22X1 OAI22X1_79 ( .A(_2030_), .B(_2471__bF_buf9), .C(_2473__bF_buf15), .D(_1964_), .Y(_1115_) );
	INVX1 INVX1_468 ( .A(micro_hash_synth_W_3__1_), .Y(_2031_) );
	OAI22X1 OAI22X1_80 ( .A(_2031_), .B(_2471__bF_buf8), .C(_2473__bF_buf14), .D(_1965_), .Y(_1116_) );
	INVX1 INVX1_469 ( .A(micro_hash_synth_W_3__2_), .Y(_2032_) );
	OAI22X1 OAI22X1_81 ( .A(_2032_), .B(_2471__bF_buf7), .C(_2473__bF_buf13), .D(_1966_), .Y(_1117_) );
	INVX1 INVX1_470 ( .A(micro_hash_synth_W_3__3_), .Y(_2033_) );
	OAI22X1 OAI22X1_82 ( .A(_2033_), .B(_2471__bF_buf6), .C(_2473__bF_buf12), .D(_1967_), .Y(_1118_) );
	INVX1 INVX1_471 ( .A(micro_hash_synth_W_3__4_), .Y(_2034_) );
	OAI22X1 OAI22X1_83 ( .A(_2034_), .B(_2471__bF_buf5), .C(_2473__bF_buf11), .D(_1968_), .Y(_1119_) );
	INVX1 INVX1_472 ( .A(micro_hash_synth_W_3__5_), .Y(_2035_) );
	OAI22X1 OAI22X1_84 ( .A(_2035_), .B(_2471__bF_buf4), .C(_2473__bF_buf10), .D(_1969_), .Y(_1120_) );
	INVX1 INVX1_473 ( .A(micro_hash_synth_W_3__6_), .Y(_2036_) );
	OAI22X1 OAI22X1_85 ( .A(_2036_), .B(_2471__bF_buf3), .C(_2473__bF_buf9), .D(_1970_), .Y(_1121_) );
	INVX1 INVX1_474 ( .A(micro_hash_synth_W_3__7_), .Y(_2037_) );
	OAI22X1 OAI22X1_86 ( .A(_2037_), .B(_2471__bF_buf2), .C(_2473__bF_buf8), .D(_1971_), .Y(_1122_) );
	INVX1 INVX1_475 ( .A(micro_hash_synth_W_4__0_), .Y(_2038_) );
	INVX1 INVX1_476 ( .A(bloque_in_32_), .Y(_2039_) );
	OAI22X1 OAI22X1_87 ( .A(_2038_), .B(_2471__bF_buf1), .C(_2473__bF_buf7), .D(_2039_), .Y(_1123_) );
	INVX1 INVX1_477 ( .A(bloque_in_33_), .Y(_2040_) );
	OAI22X1 OAI22X1_88 ( .A(_1451_), .B(_2471__bF_buf0), .C(_2473__bF_buf6), .D(_2040_), .Y(_1124_) );
	INVX1 INVX1_478 ( .A(bloque_in_34_), .Y(_2041_) );
	OAI22X1 OAI22X1_89 ( .A(_1560_), .B(_2471__bF_buf13), .C(_2473__bF_buf5), .D(_2041_), .Y(_1126_) );
	INVX1 INVX1_479 ( .A(bloque_in_35_), .Y(_2042_) );
	OAI22X1 OAI22X1_90 ( .A(_1632_), .B(_2471__bF_buf12), .C(_2473__bF_buf4), .D(_2042_), .Y(_1127_) );
	INVX1 INVX1_480 ( .A(bloque_in_36_), .Y(_2043_) );
	OAI22X1 OAI22X1_91 ( .A(_1729_), .B(_2471__bF_buf11), .C(_2473__bF_buf3), .D(_2043_), .Y(_1128_) );
	INVX1 INVX1_481 ( .A(micro_hash_synth_W_4__5_), .Y(_2044_) );
	INVX1 INVX1_482 ( .A(bloque_in_37_), .Y(_2045_) );
	OAI22X1 OAI22X1_92 ( .A(_2044_), .B(_2471__bF_buf10), .C(_2473__bF_buf2), .D(_2045_), .Y(_1129_) );
	INVX1 INVX1_483 ( .A(micro_hash_synth_W_4__6_), .Y(_2046_) );
	INVX1 INVX1_484 ( .A(bloque_in_38_), .Y(_2047_) );
	OAI22X1 OAI22X1_93 ( .A(_2046_), .B(_2471__bF_buf9), .C(_2473__bF_buf1), .D(_2047_), .Y(_1130_) );
	INVX1 INVX1_485 ( .A(micro_hash_synth_W_4__7_), .Y(_2048_) );
	INVX1 INVX1_486 ( .A(bloque_in_39_), .Y(_2049_) );
	OAI22X1 OAI22X1_94 ( .A(_2048_), .B(_2471__bF_buf8), .C(_2473__bF_buf0), .D(_2049_), .Y(_1131_) );
	INVX1 INVX1_487 ( .A(bloque_in_88_), .Y(_2050_) );
	OAI22X1 OAI22X1_95 ( .A(_2570_), .B(_2471__bF_buf7), .C(_2473__bF_buf15), .D(_2050_), .Y(_1132_) );
	INVX1 INVX1_488 ( .A(bloque_in_89_), .Y(_2051_) );
	OAI22X1 OAI22X1_96 ( .A(_2575_), .B(_2471__bF_buf6), .C(_2473__bF_buf14), .D(_2051_), .Y(_1133_) );
	INVX1 INVX1_489 ( .A(bloque_in_90_), .Y(_2052_) );
	OAI22X1 OAI22X1_97 ( .A(_2580_), .B(_2471__bF_buf5), .C(_2473__bF_buf13), .D(_2052_), .Y(_1134_) );
	INVX1 INVX1_490 ( .A(bloque_in_91_), .Y(_2053_) );
	OAI22X1 OAI22X1_98 ( .A(_2585_), .B(_2471__bF_buf4), .C(_2473__bF_buf12), .D(_2053_), .Y(_1135_) );
	INVX1 INVX1_491 ( .A(bloque_in_92_), .Y(_2054_) );
	OAI22X1 OAI22X1_99 ( .A(_2590_), .B(_2471__bF_buf3), .C(_2473__bF_buf11), .D(_2054_), .Y(_1137_) );
	INVX1 INVX1_492 ( .A(bloque_in_93_), .Y(_2055_) );
	OAI22X1 OAI22X1_100 ( .A(_2595_), .B(_2471__bF_buf2), .C(_2473__bF_buf10), .D(_2055_), .Y(_1138_) );
	INVX1 INVX1_493 ( .A(bloque_in_94_), .Y(_2056_) );
	OAI22X1 OAI22X1_101 ( .A(_2600_), .B(_2471__bF_buf1), .C(_2473__bF_buf9), .D(_2056_), .Y(_1139_) );
	INVX1 INVX1_494 ( .A(bloque_in_95_), .Y(_2057_) );
	OAI22X1 OAI22X1_102 ( .A(_2605_), .B(_2471__bF_buf0), .C(_2473__bF_buf8), .D(_2057_), .Y(_1140_) );
	INVX1 INVX1_495 ( .A(micro_hash_synth_W_10__0_), .Y(_2058_) );
	INVX1 INVX1_496 ( .A(micro_hash_synth_W_21__0_), .Y(_2059_) );
	OAI21X1 OAI21X1_523 ( .A(_2058_), .B(micro_hash_synth_W_15__0_), .C(_2059_), .Y(_2060_) );
	AOI21X1 AOI21X1_342 ( .A(_2058_), .B(micro_hash_synth_W_15__0_), .C(_2060_), .Y(_2061_) );
	OAI22X1 OAI22X1_103 ( .A(_2475_), .B(_2471__bF_buf13), .C(_2473__bF_buf7), .D(_2061_), .Y(_1141_) );
	INVX1 INVX1_497 ( .A(micro_hash_synth_W_21__1_), .Y(_2062_) );
	OAI21X1 OAI21X1_524 ( .A(_1507_), .B(micro_hash_synth_W_15__1_), .C(_2062_), .Y(_2063_) );
	AOI21X1 AOI21X1_343 ( .A(_1507_), .B(micro_hash_synth_W_15__1_), .C(_2063_), .Y(_2064_) );
	OAI22X1 OAI22X1_104 ( .A(_2480_), .B(_2471__bF_buf12), .C(_2473__bF_buf6), .D(_2064_), .Y(_1142_) );
	INVX1 INVX1_498 ( .A(micro_hash_synth_W_10__2_), .Y(_2065_) );
	INVX1 INVX1_499 ( .A(micro_hash_synth_W_21__2_), .Y(_2066_) );
	OAI21X1 OAI21X1_525 ( .A(_2065_), .B(micro_hash_synth_W_15__2_), .C(_2066_), .Y(_2067_) );
	AOI21X1 AOI21X1_344 ( .A(_2065_), .B(micro_hash_synth_W_15__2_), .C(_2067_), .Y(_2068_) );
	OAI22X1 OAI22X1_105 ( .A(_2485_), .B(_2471__bF_buf11), .C(_2473__bF_buf5), .D(_2068_), .Y(_1143_) );
	INVX1 INVX1_500 ( .A(micro_hash_synth_W_21__3_), .Y(_2069_) );
	OAI21X1 OAI21X1_526 ( .A(_1650_), .B(micro_hash_synth_W_15__3_), .C(_2069_), .Y(_2070_) );
	AOI21X1 AOI21X1_345 ( .A(_1650_), .B(micro_hash_synth_W_15__3_), .C(_2070_), .Y(_2071_) );
	OAI22X1 OAI22X1_106 ( .A(_2490_), .B(_2471__bF_buf10), .C(_2473__bF_buf4), .D(_2071_), .Y(_1144_) );
	INVX1 INVX1_501 ( .A(micro_hash_synth_W_21__4_), .Y(_2072_) );
	OAI21X1 OAI21X1_527 ( .A(_1747_), .B(micro_hash_synth_W_15__4_), .C(_2072_), .Y(_2073_) );
	AOI21X1 AOI21X1_346 ( .A(_1747_), .B(micro_hash_synth_W_15__4_), .C(_2073_), .Y(_2074_) );
	OAI22X1 OAI22X1_107 ( .A(_2495_), .B(_2471__bF_buf9), .C(_2473__bF_buf3), .D(_2074_), .Y(_1145_) );
	INVX1 INVX1_502 ( .A(micro_hash_synth_W_10__5_), .Y(_2075_) );
	INVX1 INVX1_503 ( .A(micro_hash_synth_W_21__5_), .Y(_2076_) );
	OAI21X1 OAI21X1_528 ( .A(_2075_), .B(micro_hash_synth_W_15__5_), .C(_2076_), .Y(_2077_) );
	AOI21X1 AOI21X1_347 ( .A(_2075_), .B(micro_hash_synth_W_15__5_), .C(_2077_), .Y(_2078_) );
	OAI22X1 OAI22X1_108 ( .A(_2500_), .B(_2471__bF_buf8), .C(_2473__bF_buf2), .D(_2078_), .Y(_1146_) );
	INVX1 INVX1_504 ( .A(micro_hash_synth_W_10__6_), .Y(_2079_) );
	INVX1 INVX1_505 ( .A(micro_hash_synth_W_21__6_), .Y(_2080_) );
	OAI21X1 OAI21X1_529 ( .A(_2079_), .B(micro_hash_synth_W_15__6_), .C(_2080_), .Y(_2081_) );
	AOI21X1 AOI21X1_348 ( .A(_2079_), .B(micro_hash_synth_W_15__6_), .C(_2081_), .Y(_2082_) );
	OAI22X1 OAI22X1_109 ( .A(_2505_), .B(_2471__bF_buf7), .C(_2473__bF_buf1), .D(_2082_), .Y(_1148_) );
	INVX1 INVX1_506 ( .A(micro_hash_synth_W_10__7_), .Y(_2083_) );
	INVX1 INVX1_507 ( .A(micro_hash_synth_W_21__7_), .Y(_2084_) );
	OAI21X1 OAI21X1_530 ( .A(_2083_), .B(micro_hash_synth_W_15__7_), .C(_2084_), .Y(_2085_) );
	AOI21X1 AOI21X1_349 ( .A(_2083_), .B(micro_hash_synth_W_15__7_), .C(_2085_), .Y(_2086_) );
	OAI22X1 OAI22X1_110 ( .A(_2510_), .B(_2471__bF_buf6), .C(_2473__bF_buf0), .D(_2086_), .Y(_1149_) );
	INVX1 INVX1_508 ( .A(micro_hash_synth_W_20__0_), .Y(_2087_) );
	OAI21X1 OAI21X1_531 ( .A(_2513_), .B(micro_hash_synth_W_14__0_), .C(_2087_), .Y(_2088_) );
	AOI21X1 AOI21X1_350 ( .A(_2513_), .B(micro_hash_synth_W_14__0_), .C(_2088_), .Y(_2089_) );
	OAI22X1 OAI22X1_111 ( .A(_2531_), .B(_2471__bF_buf5), .C(_2473__bF_buf15), .D(_2089_), .Y(_1150_) );
	OAI21X1 OAI21X1_532 ( .A(_2515_), .B(micro_hash_synth_W_14__1_), .C(_1424_), .Y(_2090_) );
	AOI21X1 AOI21X1_351 ( .A(_2515_), .B(micro_hash_synth_W_14__1_), .C(_2090_), .Y(_2091_) );
	OAI22X1 OAI22X1_112 ( .A(_2536_), .B(_2471__bF_buf4), .C(_2473__bF_buf14), .D(_2091_), .Y(_1151_) );
	INVX1 INVX1_509 ( .A(micro_hash_synth_W_20__2_), .Y(_2092_) );
	OAI21X1 OAI21X1_533 ( .A(_2517_), .B(micro_hash_synth_W_14__2_), .C(_2092_), .Y(_2093_) );
	AOI21X1 AOI21X1_352 ( .A(_2517_), .B(micro_hash_synth_W_14__2_), .C(_2093_), .Y(_2094_) );
	OAI22X1 OAI22X1_113 ( .A(_2541_), .B(_2471__bF_buf3), .C(_2473__bF_buf13), .D(_2094_), .Y(_1152_) );
	OAI21X1 OAI21X1_534 ( .A(_2519_), .B(micro_hash_synth_W_14__3_), .C(_1603_), .Y(_2095_) );
	AOI21X1 AOI21X1_353 ( .A(_2519_), .B(micro_hash_synth_W_14__3_), .C(_2095_), .Y(_2096_) );
	OAI22X1 OAI22X1_114 ( .A(_2546_), .B(_2471__bF_buf2), .C(_2473__bF_buf12), .D(_2096_), .Y(_1153_) );
	OAI21X1 OAI21X1_535 ( .A(_2521_), .B(micro_hash_synth_W_14__4_), .C(_1706_), .Y(_2097_) );
	AOI21X1 AOI21X1_354 ( .A(_2521_), .B(micro_hash_synth_W_14__4_), .C(_2097_), .Y(_2098_) );
	OAI22X1 OAI22X1_115 ( .A(_2551_), .B(_2471__bF_buf1), .C(_2473__bF_buf11), .D(_2098_), .Y(_1154_) );
	INVX1 INVX1_510 ( .A(micro_hash_synth_W_20__5_), .Y(_2099_) );
	OAI21X1 OAI21X1_536 ( .A(_2523_), .B(micro_hash_synth_W_14__5_), .C(_2099_), .Y(_2100_) );
	AOI21X1 AOI21X1_355 ( .A(_2523_), .B(micro_hash_synth_W_14__5_), .C(_2100_), .Y(_2101_) );
	OAI22X1 OAI22X1_116 ( .A(_2556_), .B(_2471__bF_buf0), .C(_2473__bF_buf10), .D(_2101_), .Y(_1155_) );
	INVX1 INVX1_511 ( .A(micro_hash_synth_W_20__6_), .Y(_2102_) );
	OAI21X1 OAI21X1_537 ( .A(_2525_), .B(micro_hash_synth_W_14__6_), .C(_2102_), .Y(_2103_) );
	AOI21X1 AOI21X1_356 ( .A(_2525_), .B(micro_hash_synth_W_14__6_), .C(_2103_), .Y(_2104_) );
	OAI22X1 OAI22X1_117 ( .A(_2561_), .B(_2471__bF_buf13), .C(_2473__bF_buf9), .D(_2104_), .Y(_1156_) );
	INVX1 INVX1_512 ( .A(micro_hash_synth_W_20__7_), .Y(_2105_) );
	OAI21X1 OAI21X1_538 ( .A(_2527_), .B(micro_hash_synth_W_14__7_), .C(_2105_), .Y(_2106_) );
	AOI21X1 AOI21X1_357 ( .A(_2527_), .B(micro_hash_synth_W_14__7_), .C(_2106_), .Y(_2107_) );
	OAI22X1 OAI22X1_118 ( .A(_2566_), .B(_2471__bF_buf12), .C(_2473__bF_buf8), .D(_2107_), .Y(_1157_) );
	INVX1 INVX1_513 ( .A(micro_hash_synth_W_8__0_), .Y(_2108_) );
	INVX1 INVX1_514 ( .A(bloque_in_64_), .Y(_2109_) );
	OAI22X1 OAI22X1_119 ( .A(_2108_), .B(_2471__bF_buf11), .C(_2473__bF_buf7), .D(_2109_), .Y(_1159_) );
	INVX1 INVX1_515 ( .A(bloque_in_65_), .Y(_2110_) );
	OAI22X1 OAI22X1_120 ( .A(_1464_), .B(_2471__bF_buf10), .C(_2473__bF_buf6), .D(_2110_), .Y(_1160_) );
	INVX1 INVX1_516 ( .A(micro_hash_synth_W_8__2_), .Y(_2111_) );
	INVX1 INVX1_517 ( .A(bloque_in_66_), .Y(_2112_) );
	OAI22X1 OAI22X1_121 ( .A(_2111_), .B(_2471__bF_buf9), .C(_2473__bF_buf5), .D(_2112_), .Y(_1161_) );
	INVX1 INVX1_518 ( .A(bloque_in_67_), .Y(_2113_) );
	OAI22X1 OAI22X1_122 ( .A(_1653_), .B(_2471__bF_buf8), .C(_2473__bF_buf4), .D(_2113_), .Y(_1162_) );
	INVX1 INVX1_519 ( .A(bloque_in_68_), .Y(_2114_) );
	OAI22X1 OAI22X1_123 ( .A(_1750_), .B(_2471__bF_buf7), .C(_2473__bF_buf3), .D(_2114_), .Y(_1163_) );
	INVX1 INVX1_520 ( .A(micro_hash_synth_W_8__5_), .Y(_2115_) );
	INVX1 INVX1_521 ( .A(bloque_in_69_), .Y(_2116_) );
	OAI22X1 OAI22X1_124 ( .A(_2115_), .B(_2471__bF_buf6), .C(_2473__bF_buf2), .D(_2116_), .Y(_1164_) );
	INVX1 INVX1_522 ( .A(micro_hash_synth_W_8__6_), .Y(_2117_) );
	INVX1 INVX1_523 ( .A(bloque_in_70_), .Y(_2118_) );
	OAI22X1 OAI22X1_125 ( .A(_2117_), .B(_2471__bF_buf5), .C(_2473__bF_buf1), .D(_2118_), .Y(_1165_) );
	INVX1 INVX1_524 ( .A(micro_hash_synth_W_8__7_), .Y(_2119_) );
	INVX1 INVX1_525 ( .A(bloque_in_71_), .Y(_2120_) );
	OAI22X1 OAI22X1_126 ( .A(_2119_), .B(_2471__bF_buf4), .C(_2473__bF_buf0), .D(_2120_), .Y(_1166_) );
	INVX1 INVX1_526 ( .A(micro_hash_synth_W_19__0_), .Y(_2121_) );
	OAI21X1 OAI21X1_539 ( .A(_2108_), .B(micro_hash_synth_W_13__0_), .C(_2121_), .Y(_2122_) );
	AOI21X1 AOI21X1_358 ( .A(micro_hash_synth_W_13__0_), .B(_2108_), .C(_2122_), .Y(_2123_) );
	OAI22X1 OAI22X1_127 ( .A(_2571_), .B(_2471__bF_buf3), .C(_2473__bF_buf15), .D(_2123_), .Y(_1167_) );
	INVX1 INVX1_527 ( .A(micro_hash_synth_W_19__1_), .Y(_2124_) );
	OAI21X1 OAI21X1_540 ( .A(_1464_), .B(micro_hash_synth_W_13__1_), .C(_2124_), .Y(_2125_) );
	AOI21X1 AOI21X1_359 ( .A(micro_hash_synth_W_13__1_), .B(_1464_), .C(_2125_), .Y(_2126_) );
	OAI22X1 OAI22X1_128 ( .A(_2576_), .B(_2471__bF_buf2), .C(_2473__bF_buf14), .D(_2126_), .Y(_1168_) );
	INVX1 INVX1_528 ( .A(micro_hash_synth_W_19__2_), .Y(_2127_) );
	OAI21X1 OAI21X1_541 ( .A(_2111_), .B(micro_hash_synth_W_13__2_), .C(_2127_), .Y(_2128_) );
	AOI21X1 AOI21X1_360 ( .A(micro_hash_synth_W_13__2_), .B(_2111_), .C(_2128_), .Y(_2129_) );
	OAI22X1 OAI22X1_129 ( .A(_2581_), .B(_2471__bF_buf1), .C(_2473__bF_buf13), .D(_2129_), .Y(_1170_) );
	INVX1 INVX1_529 ( .A(micro_hash_synth_W_19__3_), .Y(_2130_) );
	OAI21X1 OAI21X1_542 ( .A(_1653_), .B(micro_hash_synth_W_13__3_), .C(_2130_), .Y(_2131_) );
	AOI21X1 AOI21X1_361 ( .A(micro_hash_synth_W_13__3_), .B(_1653_), .C(_2131_), .Y(_2132_) );
	OAI22X1 OAI22X1_130 ( .A(_2586_), .B(_2471__bF_buf0), .C(_2473__bF_buf12), .D(_2132_), .Y(_1171_) );
	INVX1 INVX1_530 ( .A(micro_hash_synth_W_19__4_), .Y(_2133_) );
	OAI21X1 OAI21X1_543 ( .A(_1750_), .B(micro_hash_synth_W_13__4_), .C(_2133_), .Y(_2134_) );
	AOI21X1 AOI21X1_362 ( .A(micro_hash_synth_W_13__4_), .B(_1750_), .C(_2134_), .Y(_2135_) );
	OAI22X1 OAI22X1_131 ( .A(_2591_), .B(_2471__bF_buf13), .C(_2473__bF_buf11), .D(_2135_), .Y(_1172_) );
	INVX1 INVX1_531 ( .A(micro_hash_synth_W_19__5_), .Y(_2136_) );
	OAI21X1 OAI21X1_544 ( .A(_2115_), .B(micro_hash_synth_W_13__5_), .C(_2136_), .Y(_2137_) );
	AOI21X1 AOI21X1_363 ( .A(micro_hash_synth_W_13__5_), .B(_2115_), .C(_2137_), .Y(_2138_) );
	OAI22X1 OAI22X1_132 ( .A(_2596_), .B(_2471__bF_buf12), .C(_2473__bF_buf10), .D(_2138_), .Y(_1173_) );
	INVX1 INVX1_532 ( .A(micro_hash_synth_W_19__6_), .Y(_2139_) );
	OAI21X1 OAI21X1_545 ( .A(_2117_), .B(micro_hash_synth_W_13__6_), .C(_2139_), .Y(_2140_) );
	AOI21X1 AOI21X1_364 ( .A(micro_hash_synth_W_13__6_), .B(_2117_), .C(_2140_), .Y(_2141_) );
	OAI22X1 OAI22X1_133 ( .A(_2601_), .B(_2471__bF_buf11), .C(_2473__bF_buf9), .D(_2141_), .Y(_1174_) );
	INVX1 INVX1_533 ( .A(micro_hash_synth_W_19__7_), .Y(_2142_) );
	OAI21X1 OAI21X1_546 ( .A(_2119_), .B(micro_hash_synth_W_13__7_), .C(_2142_), .Y(_2143_) );
	AOI21X1 AOI21X1_365 ( .A(micro_hash_synth_W_13__7_), .B(_2119_), .C(_2143_), .Y(_2144_) );
	OAI22X1 OAI22X1_134 ( .A(_2606_), .B(_2471__bF_buf10), .C(_2473__bF_buf8), .D(_2144_), .Y(_1175_) );
	INVX1 INVX1_534 ( .A(micro_hash_synth_W_5__0_), .Y(_2145_) );
	INVX1 INVX1_535 ( .A(bloque_in_40_), .Y(_2146_) );
	OAI22X1 OAI22X1_135 ( .A(_2145_), .B(_2471__bF_buf9), .C(_2473__bF_buf7), .D(_2146_), .Y(_1181_) );
	INVX1 INVX1_536 ( .A(bloque_in_41_), .Y(_2147_) );
	OAI22X1 OAI22X1_136 ( .A(_1453_), .B(_2471__bF_buf8), .C(_2473__bF_buf6), .D(_2147_), .Y(_1182_) );
	INVX1 INVX1_537 ( .A(micro_hash_synth_W_5__2_), .Y(_2148_) );
	INVX1 INVX1_538 ( .A(bloque_in_42_), .Y(_2149_) );
	OAI22X1 OAI22X1_137 ( .A(_2148_), .B(_2471__bF_buf7), .C(_2473__bF_buf5), .D(_2149_), .Y(_1183_) );
	INVX1 INVX1_539 ( .A(micro_hash_synth_W_5__3_), .Y(_2150_) );
	INVX1 INVX1_540 ( .A(bloque_in_43_), .Y(_2151_) );
	OAI22X1 OAI22X1_138 ( .A(_2150_), .B(_2471__bF_buf6), .C(_2473__bF_buf4), .D(_2151_), .Y(_1184_) );
	INVX1 INVX1_541 ( .A(micro_hash_synth_W_5__4_), .Y(_2152_) );
	INVX1 INVX1_542 ( .A(bloque_in_44_), .Y(_2153_) );
	OAI22X1 OAI22X1_139 ( .A(_2152_), .B(_2471__bF_buf5), .C(_2473__bF_buf3), .D(_2153_), .Y(_1185_) );
	INVX1 INVX1_543 ( .A(micro_hash_synth_W_5__5_), .Y(_2154_) );
	INVX1 INVX1_544 ( .A(bloque_in_45_), .Y(_2155_) );
	OAI22X1 OAI22X1_140 ( .A(_2154_), .B(_2471__bF_buf4), .C(_2473__bF_buf2), .D(_2155_), .Y(_1186_) );
	INVX1 INVX1_545 ( .A(micro_hash_synth_W_5__6_), .Y(_2156_) );
	INVX1 INVX1_546 ( .A(bloque_in_46_), .Y(_2157_) );
	OAI22X1 OAI22X1_141 ( .A(_2156_), .B(_2471__bF_buf3), .C(_2473__bF_buf1), .D(_2157_), .Y(_1187_) );
	INVX1 INVX1_547 ( .A(micro_hash_synth_W_5__7_), .Y(_2158_) );
	INVX1 INVX1_548 ( .A(bloque_in_47_), .Y(_2159_) );
	OAI22X1 OAI22X1_142 ( .A(_2158_), .B(_2471__bF_buf2), .C(_2473__bF_buf0), .D(_2159_), .Y(_1189_) );
	INVX1 INVX1_549 ( .A(micro_hash_synth_W_7__0_), .Y(_2160_) );
	INVX1 INVX1_550 ( .A(micro_hash_synth_W_18__0_), .Y(_2161_) );
	OAI21X1 OAI21X1_547 ( .A(_2160_), .B(micro_hash_synth_W_12__0_), .C(_2161_), .Y(_2162_) );
	AOI21X1 AOI21X1_366 ( .A(micro_hash_synth_W_12__0_), .B(_2160_), .C(_2162_), .Y(_2163_) );
	OAI22X1 OAI22X1_143 ( .A(_2059_), .B(_2471__bF_buf1), .C(_2473__bF_buf15), .D(_2163_), .Y(_942_) );
	INVX1 INVX1_551 ( .A(micro_hash_synth_W_7__1_), .Y(_2164_) );
	OAI21X1 OAI21X1_548 ( .A(_2164_), .B(micro_hash_synth_W_12__1_), .C(_1473_), .Y(_2165_) );
	AOI21X1 AOI21X1_367 ( .A(micro_hash_synth_W_12__1_), .B(_2164_), .C(_2165_), .Y(_2166_) );
	OAI22X1 OAI22X1_144 ( .A(_2062_), .B(_2471__bF_buf0), .C(_2473__bF_buf14), .D(_2166_), .Y(_943_) );
	INVX1 INVX1_552 ( .A(micro_hash_synth_W_7__2_), .Y(_2167_) );
	INVX1 INVX1_553 ( .A(micro_hash_synth_W_18__2_), .Y(_2168_) );
	OAI21X1 OAI21X1_549 ( .A(_2167_), .B(micro_hash_synth_W_12__2_), .C(_2168_), .Y(_2169_) );
	AOI21X1 AOI21X1_368 ( .A(micro_hash_synth_W_12__2_), .B(_2167_), .C(_2169_), .Y(_2170_) );
	OAI22X1 OAI22X1_145 ( .A(_2066_), .B(_2471__bF_buf13), .C(_2473__bF_buf13), .D(_2170_), .Y(_944_) );
	INVX1 INVX1_554 ( .A(micro_hash_synth_W_7__3_), .Y(_2171_) );
	OAI21X1 OAI21X1_550 ( .A(_2171_), .B(micro_hash_synth_W_12__3_), .C(_1607_), .Y(_2172_) );
	AOI21X1 AOI21X1_369 ( .A(micro_hash_synth_W_12__3_), .B(_2171_), .C(_2172_), .Y(_2173_) );
	OAI22X1 OAI22X1_146 ( .A(_2069_), .B(_2471__bF_buf12), .C(_2473__bF_buf12), .D(_2173_), .Y(_945_) );
	INVX1 INVX1_555 ( .A(micro_hash_synth_W_7__4_), .Y(_2174_) );
	OAI21X1 OAI21X1_551 ( .A(_2174_), .B(micro_hash_synth_W_12__4_), .C(_1700_), .Y(_2175_) );
	AOI21X1 AOI21X1_370 ( .A(micro_hash_synth_W_12__4_), .B(_2174_), .C(_2175_), .Y(_2176_) );
	OAI22X1 OAI22X1_147 ( .A(_2072_), .B(_2471__bF_buf11), .C(_2473__bF_buf11), .D(_2176_), .Y(_946_) );
	INVX1 INVX1_556 ( .A(micro_hash_synth_W_7__5_), .Y(_2177_) );
	INVX1 INVX1_557 ( .A(micro_hash_synth_W_18__5_), .Y(_2178_) );
	OAI21X1 OAI21X1_552 ( .A(_2177_), .B(micro_hash_synth_W_12__5_), .C(_2178_), .Y(_2179_) );
	AOI21X1 AOI21X1_371 ( .A(micro_hash_synth_W_12__5_), .B(_2177_), .C(_2179_), .Y(_2180_) );
	OAI22X1 OAI22X1_148 ( .A(_2076_), .B(_2471__bF_buf10), .C(_2473__bF_buf10), .D(_2180_), .Y(_947_) );
	INVX1 INVX1_558 ( .A(micro_hash_synth_W_7__6_), .Y(_2181_) );
	INVX1 INVX1_559 ( .A(micro_hash_synth_W_18__6_), .Y(_2182_) );
	OAI21X1 OAI21X1_553 ( .A(_2181_), .B(micro_hash_synth_W_12__6_), .C(_2182_), .Y(_2183_) );
	AOI21X1 AOI21X1_372 ( .A(micro_hash_synth_W_12__6_), .B(_2181_), .C(_2183_), .Y(_2184_) );
	OAI22X1 OAI22X1_149 ( .A(_2080_), .B(_2471__bF_buf9), .C(_2473__bF_buf9), .D(_2184_), .Y(_948_) );
	INVX1 INVX1_560 ( .A(micro_hash_synth_W_7__7_), .Y(_2185_) );
	INVX1 INVX1_561 ( .A(micro_hash_synth_W_18__7_), .Y(_2186_) );
	OAI21X1 OAI21X1_554 ( .A(_2185_), .B(micro_hash_synth_W_12__7_), .C(_2186_), .Y(_2187_) );
	AOI21X1 AOI21X1_373 ( .A(micro_hash_synth_W_12__7_), .B(_2185_), .C(_2187_), .Y(_2188_) );
	OAI22X1 OAI22X1_150 ( .A(_2084_), .B(_2471__bF_buf8), .C(_2473__bF_buf8), .D(_2188_), .Y(_949_) );
	INVX8 INVX8_4 ( .A(_2471__bF_buf7), .Y(_2189_) );
	NAND2X1 NAND2X1_230 ( .A(micro_hash_synth_W_0__0_), .B(_2189__bF_buf4), .Y(_2190_) );
	OAI21X1 OAI21X1_555 ( .A(_1940_), .B(_2473__bF_buf7), .C(_2190_), .Y(_951_) );
	OAI22X1 OAI22X1_151 ( .A(_1493_), .B(_2471__bF_buf6), .C(_2473__bF_buf6), .D(_1941_), .Y(_952_) );
	NAND2X1 NAND2X1_231 ( .A(micro_hash_synth_W_0__2_), .B(_2189__bF_buf3), .Y(_2191_) );
	OAI21X1 OAI21X1_556 ( .A(_1942_), .B(_2473__bF_buf5), .C(_2191_), .Y(_953_) );
	OAI22X1 OAI22X1_152 ( .A(_1639_), .B(_2471__bF_buf5), .C(_2473__bF_buf4), .D(_1943_), .Y(_954_) );
	OAI22X1 OAI22X1_153 ( .A(_1736_), .B(_2471__bF_buf4), .C(_2473__bF_buf3), .D(_1944_), .Y(_956_) );
	NAND2X1 NAND2X1_232 ( .A(micro_hash_synth_W_0__5_), .B(_2189__bF_buf2), .Y(_2192_) );
	OAI21X1 OAI21X1_557 ( .A(_1945_), .B(_2473__bF_buf2), .C(_2192_), .Y(_957_) );
	NAND2X1 NAND2X1_233 ( .A(micro_hash_synth_W_0__6_), .B(_2189__bF_buf1), .Y(_2193_) );
	OAI21X1 OAI21X1_558 ( .A(_1946_), .B(_2473__bF_buf1), .C(_2193_), .Y(_958_) );
	NAND2X1 NAND2X1_234 ( .A(micro_hash_synth_W_0__7_), .B(_2189__bF_buf0), .Y(_2194_) );
	OAI21X1 OAI21X1_559 ( .A(_1947_), .B(_2473__bF_buf0), .C(_2194_), .Y(_959_) );
	INVX1 INVX1_562 ( .A(micro_hash_synth_W_6__0_), .Y(_2195_) );
	INVX1 INVX1_563 ( .A(micro_hash_synth_W_17__0_), .Y(_2196_) );
	OAI21X1 OAI21X1_560 ( .A(_2195_), .B(micro_hash_synth_W_11__0_), .C(_2196_), .Y(_2197_) );
	AOI21X1 AOI21X1_374 ( .A(micro_hash_synth_W_11__0_), .B(_2195_), .C(_2197_), .Y(_2198_) );
	OAI22X1 OAI22X1_154 ( .A(_2087_), .B(_2471__bF_buf3), .C(_2473__bF_buf15), .D(_2198_), .Y(_960_) );
	OAI21X1 OAI21X1_561 ( .A(_1487_), .B(micro_hash_synth_W_11__1_), .C(_1432_), .Y(_2199_) );
	AOI21X1 AOI21X1_375 ( .A(micro_hash_synth_W_11__1_), .B(_1487_), .C(_2199_), .Y(_2200_) );
	OAI22X1 OAI22X1_155 ( .A(_1424_), .B(_2471__bF_buf2), .C(_2473__bF_buf14), .D(_2200_), .Y(_961_) );
	OAI21X1 OAI21X1_562 ( .A(_1557_), .B(micro_hash_synth_W_11__2_), .C(_1529_), .Y(_2201_) );
	AOI21X1 AOI21X1_376 ( .A(micro_hash_synth_W_11__2_), .B(_1557_), .C(_2201_), .Y(_2202_) );
	OAI22X1 OAI22X1_156 ( .A(_2092_), .B(_2471__bF_buf1), .C(_2473__bF_buf13), .D(_2202_), .Y(_962_) );
	INVX1 INVX1_564 ( .A(micro_hash_synth_W_17__3_), .Y(_2203_) );
	OAI21X1 OAI21X1_563 ( .A(_1629_), .B(micro_hash_synth_W_11__3_), .C(_2203_), .Y(_2204_) );
	AOI21X1 AOI21X1_377 ( .A(micro_hash_synth_W_11__3_), .B(_1629_), .C(_2204_), .Y(_2205_) );
	OAI22X1 OAI22X1_157 ( .A(_1603_), .B(_2471__bF_buf0), .C(_2473__bF_buf12), .D(_2205_), .Y(_963_) );
	INVX1 INVX1_565 ( .A(micro_hash_synth_W_17__4_), .Y(_2206_) );
	OAI21X1 OAI21X1_564 ( .A(_1726_), .B(micro_hash_synth_W_11__4_), .C(_2206_), .Y(_2207_) );
	AOI21X1 AOI21X1_378 ( .A(micro_hash_synth_W_11__4_), .B(_1726_), .C(_2207_), .Y(_2208_) );
	OAI22X1 OAI22X1_158 ( .A(_1706_), .B(_2471__bF_buf13), .C(_2473__bF_buf11), .D(_2208_), .Y(_964_) );
	INVX1 INVX1_566 ( .A(micro_hash_synth_W_6__5_), .Y(_2209_) );
	INVX1 INVX1_567 ( .A(micro_hash_synth_W_17__5_), .Y(_2210_) );
	OAI21X1 OAI21X1_565 ( .A(_2209_), .B(micro_hash_synth_W_11__5_), .C(_2210_), .Y(_2211_) );
	AOI21X1 AOI21X1_379 ( .A(micro_hash_synth_W_11__5_), .B(_2209_), .C(_2211_), .Y(_2212_) );
	OAI22X1 OAI22X1_159 ( .A(_2099_), .B(_2471__bF_buf12), .C(_2473__bF_buf10), .D(_2212_), .Y(_965_) );
	INVX1 INVX1_568 ( .A(micro_hash_synth_W_6__6_), .Y(_2213_) );
	INVX1 INVX1_569 ( .A(micro_hash_synth_W_17__6_), .Y(_2214_) );
	OAI21X1 OAI21X1_566 ( .A(_2213_), .B(micro_hash_synth_W_11__6_), .C(_2214_), .Y(_2215_) );
	AOI21X1 AOI21X1_380 ( .A(micro_hash_synth_W_11__6_), .B(_2213_), .C(_2215_), .Y(_2216_) );
	OAI22X1 OAI22X1_160 ( .A(_2102_), .B(_2471__bF_buf11), .C(_2473__bF_buf9), .D(_2216_), .Y(_966_) );
	INVX1 INVX1_570 ( .A(micro_hash_synth_W_6__7_), .Y(_2217_) );
	INVX1 INVX1_571 ( .A(micro_hash_synth_W_17__7_), .Y(_2218_) );
	OAI21X1 OAI21X1_567 ( .A(_2217_), .B(micro_hash_synth_W_11__7_), .C(_2218_), .Y(_2219_) );
	AOI21X1 AOI21X1_381 ( .A(micro_hash_synth_W_11__7_), .B(_2217_), .C(_2219_), .Y(_2220_) );
	OAI22X1 OAI22X1_161 ( .A(_2105_), .B(_2471__bF_buf10), .C(_2473__bF_buf8), .D(_2220_), .Y(_967_) );
	INVX1 INVX1_572 ( .A(bloque_in_48_), .Y(_2221_) );
	OAI22X1 OAI22X1_162 ( .A(_2195_), .B(_2471__bF_buf9), .C(_2473__bF_buf7), .D(_2221_), .Y(_968_) );
	INVX1 INVX1_573 ( .A(bloque_in_49_), .Y(_2222_) );
	OAI22X1 OAI22X1_163 ( .A(_1487_), .B(_2471__bF_buf8), .C(_2473__bF_buf6), .D(_2222_), .Y(_969_) );
	INVX1 INVX1_574 ( .A(bloque_in_50_), .Y(_2223_) );
	OAI22X1 OAI22X1_164 ( .A(_1557_), .B(_2471__bF_buf7), .C(_2473__bF_buf5), .D(_2223_), .Y(_970_) );
	INVX1 INVX1_575 ( .A(bloque_in_51_), .Y(_2224_) );
	OAI22X1 OAI22X1_165 ( .A(_1629_), .B(_2471__bF_buf6), .C(_2473__bF_buf4), .D(_2224_), .Y(_972_) );
	INVX1 INVX1_576 ( .A(bloque_in_52_), .Y(_2225_) );
	OAI22X1 OAI22X1_166 ( .A(_1726_), .B(_2471__bF_buf5), .C(_2473__bF_buf3), .D(_2225_), .Y(_973_) );
	INVX1 INVX1_577 ( .A(bloque_in_53_), .Y(_2226_) );
	OAI22X1 OAI22X1_167 ( .A(_2209_), .B(_2471__bF_buf4), .C(_2473__bF_buf2), .D(_2226_), .Y(_974_) );
	INVX1 INVX1_578 ( .A(bloque_in_54_), .Y(_2227_) );
	OAI22X1 OAI22X1_168 ( .A(_2213_), .B(_2471__bF_buf3), .C(_2473__bF_buf1), .D(_2227_), .Y(_975_) );
	INVX1 INVX1_579 ( .A(bloque_in_55_), .Y(_2228_) );
	OAI22X1 OAI22X1_169 ( .A(_2217_), .B(_2471__bF_buf2), .C(_2473__bF_buf0), .D(_2228_), .Y(_976_) );
	INVX1 INVX1_580 ( .A(micro_hash_synth_W_15__0_), .Y(_2229_) );
	INVX1 INVX1_581 ( .A(bloque_in_120_), .Y(_2230_) );
	OAI22X1 OAI22X1_170 ( .A(_2229_), .B(_2471__bF_buf1), .C(_2473__bF_buf15), .D(_2230_), .Y(_977_) );
	INVX1 INVX1_582 ( .A(micro_hash_synth_W_15__1_), .Y(_2231_) );
	INVX1 INVX1_583 ( .A(bloque_in_121_), .Y(_2232_) );
	OAI22X1 OAI22X1_171 ( .A(_2231_), .B(_2471__bF_buf0), .C(_2473__bF_buf14), .D(_2232_), .Y(_978_) );
	INVX1 INVX1_584 ( .A(micro_hash_synth_W_15__2_), .Y(_2233_) );
	INVX1 INVX1_585 ( .A(bloque_in_122_), .Y(_2234_) );
	OAI22X1 OAI22X1_172 ( .A(_2233_), .B(_2471__bF_buf13), .C(_2473__bF_buf13), .D(_2234_), .Y(_979_) );
	INVX1 INVX1_586 ( .A(micro_hash_synth_W_15__3_), .Y(_2235_) );
	INVX1 INVX1_587 ( .A(bloque_in_123_), .Y(_2236_) );
	OAI22X1 OAI22X1_173 ( .A(_2235_), .B(_2471__bF_buf12), .C(_2473__bF_buf12), .D(_2236_), .Y(_980_) );
	INVX1 INVX1_588 ( .A(micro_hash_synth_W_15__4_), .Y(_2237_) );
	INVX1 INVX1_589 ( .A(bloque_in_124_), .Y(_2238_) );
	OAI22X1 OAI22X1_174 ( .A(_2237_), .B(_2471__bF_buf11), .C(_2473__bF_buf11), .D(_2238_), .Y(_981_) );
	INVX1 INVX1_590 ( .A(micro_hash_synth_W_15__5_), .Y(_2239_) );
	INVX1 INVX1_591 ( .A(bloque_in_125_), .Y(_2240_) );
	OAI22X1 OAI22X1_175 ( .A(_2239_), .B(_2471__bF_buf10), .C(_2473__bF_buf10), .D(_2240_), .Y(_982_) );
	INVX1 INVX1_592 ( .A(micro_hash_synth_W_15__6_), .Y(_2241_) );
	INVX1 INVX1_593 ( .A(bloque_in_126_), .Y(_2242_) );
	OAI22X1 OAI22X1_176 ( .A(_2241_), .B(_2471__bF_buf9), .C(_2473__bF_buf9), .D(_2242_), .Y(_983_) );
	INVX1 INVX1_594 ( .A(micro_hash_synth_W_15__7_), .Y(_2243_) );
	INVX1 INVX1_595 ( .A(bloque_in_127_), .Y(_2244_) );
	OAI22X1 OAI22X1_177 ( .A(_2243_), .B(_2471__bF_buf8), .C(_2473__bF_buf8), .D(_2244_), .Y(_984_) );
	INVX1 INVX1_596 ( .A(micro_hash_synth_W_16__0_), .Y(_2245_) );
	OAI21X1 OAI21X1_568 ( .A(_2145_), .B(micro_hash_synth_W_10__0_), .C(_2245_), .Y(_2246_) );
	AOI21X1 AOI21X1_382 ( .A(_2145_), .B(micro_hash_synth_W_10__0_), .C(_2246_), .Y(_2247_) );
	OAI22X1 OAI22X1_178 ( .A(_2121_), .B(_2471__bF_buf7), .C(_2473__bF_buf7), .D(_2247_), .Y(_985_) );
	OAI21X1 OAI21X1_569 ( .A(_1453_), .B(micro_hash_synth_W_10__1_), .C(_1429_), .Y(_2248_) );
	AOI21X1 AOI21X1_383 ( .A(_1453_), .B(micro_hash_synth_W_10__1_), .C(_2248_), .Y(_2249_) );
	OAI22X1 OAI22X1_179 ( .A(_2124_), .B(_2471__bF_buf6), .C(_2473__bF_buf6), .D(_2249_), .Y(_986_) );
	OAI21X1 OAI21X1_570 ( .A(_2148_), .B(micro_hash_synth_W_10__2_), .C(_1527_), .Y(_2250_) );
	AOI21X1 AOI21X1_384 ( .A(_2148_), .B(micro_hash_synth_W_10__2_), .C(_2250_), .Y(_2251_) );
	OAI22X1 OAI22X1_180 ( .A(_2127_), .B(_2471__bF_buf5), .C(_2473__bF_buf5), .D(_2251_), .Y(_988_) );
	OAI21X1 OAI21X1_571 ( .A(_2150_), .B(micro_hash_synth_W_10__3_), .C(_1610_), .Y(_2252_) );
	AOI21X1 AOI21X1_385 ( .A(_2150_), .B(micro_hash_synth_W_10__3_), .C(_2252_), .Y(_2253_) );
	OAI22X1 OAI22X1_181 ( .A(_2130_), .B(_2471__bF_buf4), .C(_2473__bF_buf4), .D(_2253_), .Y(_989_) );
	OAI21X1 OAI21X1_572 ( .A(_2152_), .B(micro_hash_synth_W_10__4_), .C(_1697_), .Y(_2254_) );
	AOI21X1 AOI21X1_386 ( .A(_2152_), .B(micro_hash_synth_W_10__4_), .C(_2254_), .Y(_2255_) );
	OAI22X1 OAI22X1_182 ( .A(_2133_), .B(_2471__bF_buf3), .C(_2473__bF_buf3), .D(_2255_), .Y(_990_) );
	INVX1 INVX1_597 ( .A(micro_hash_synth_W_16__5_), .Y(_2256_) );
	OAI21X1 OAI21X1_573 ( .A(_2154_), .B(micro_hash_synth_W_10__5_), .C(_2256_), .Y(_2257_) );
	AOI21X1 AOI21X1_387 ( .A(_2154_), .B(micro_hash_synth_W_10__5_), .C(_2257_), .Y(_2258_) );
	OAI22X1 OAI22X1_183 ( .A(_2136_), .B(_2471__bF_buf2), .C(_2473__bF_buf2), .D(_2258_), .Y(_991_) );
	INVX1 INVX1_598 ( .A(micro_hash_synth_W_16__6_), .Y(_2259_) );
	OAI21X1 OAI21X1_574 ( .A(_2156_), .B(micro_hash_synth_W_10__6_), .C(_2259_), .Y(_2260_) );
	AOI21X1 AOI21X1_388 ( .A(_2156_), .B(micro_hash_synth_W_10__6_), .C(_2260_), .Y(_2261_) );
	OAI22X1 OAI22X1_184 ( .A(_2139_), .B(_2471__bF_buf1), .C(_2473__bF_buf1), .D(_2261_), .Y(_992_) );
	INVX1 INVX1_599 ( .A(micro_hash_synth_W_16__7_), .Y(_2262_) );
	OAI21X1 OAI21X1_575 ( .A(_2158_), .B(micro_hash_synth_W_10__7_), .C(_2262_), .Y(_2263_) );
	AOI21X1 AOI21X1_389 ( .A(_2158_), .B(micro_hash_synth_W_10__7_), .C(_2263_), .Y(_2264_) );
	OAI22X1 OAI22X1_185 ( .A(_2142_), .B(_2471__bF_buf0), .C(_2473__bF_buf0), .D(_2264_), .Y(_993_) );
	NAND2X1 NAND2X1_235 ( .A(micro_hash_synth_W_1__0_), .B(_2189__bF_buf4), .Y(_2265_) );
	OAI21X1 OAI21X1_576 ( .A(_1948_), .B(_2473__bF_buf15), .C(_2265_), .Y(_994_) );
	NAND2X1 NAND2X1_236 ( .A(micro_hash_synth_W_1__1_), .B(_2189__bF_buf3), .Y(_2266_) );
	OAI21X1 OAI21X1_577 ( .A(_1949_), .B(_2473__bF_buf14), .C(_2266_), .Y(_995_) );
	NAND2X1 NAND2X1_237 ( .A(micro_hash_synth_W_1__2_), .B(_2189__bF_buf2), .Y(_2267_) );
	OAI21X1 OAI21X1_578 ( .A(_1950_), .B(_2473__bF_buf13), .C(_2267_), .Y(_996_) );
	NAND2X1 NAND2X1_238 ( .A(micro_hash_synth_W_1__3_), .B(_2189__bF_buf1), .Y(_2268_) );
	OAI21X1 OAI21X1_579 ( .A(_1951_), .B(_2473__bF_buf12), .C(_2268_), .Y(_997_) );
	NAND2X1 NAND2X1_239 ( .A(micro_hash_synth_W_1__4_), .B(_2189__bF_buf0), .Y(_2269_) );
	OAI21X1 OAI21X1_580 ( .A(_1952_), .B(_2473__bF_buf11), .C(_2269_), .Y(_998_) );
	NAND2X1 NAND2X1_240 ( .A(micro_hash_synth_W_1__5_), .B(_2189__bF_buf4), .Y(_2270_) );
	OAI21X1 OAI21X1_581 ( .A(_1953_), .B(_2473__bF_buf10), .C(_2270_), .Y(_999_) );
	NAND2X1 NAND2X1_241 ( .A(micro_hash_synth_W_1__6_), .B(_2189__bF_buf3), .Y(_2271_) );
	OAI21X1 OAI21X1_582 ( .A(_1954_), .B(_2473__bF_buf9), .C(_2271_), .Y(_1000_) );
	NAND2X1 NAND2X1_242 ( .A(micro_hash_synth_W_1__7_), .B(_2189__bF_buf2), .Y(_2272_) );
	OAI21X1 OAI21X1_583 ( .A(_1955_), .B(_2473__bF_buf8), .C(_2272_), .Y(_1001_) );
	OAI21X1 OAI21X1_584 ( .A(_2038_), .B(micro_hash_synth_W_9__0_), .C(_2229_), .Y(_2273_) );
	AOI21X1 AOI21X1_390 ( .A(micro_hash_synth_W_9__0_), .B(_2038_), .C(_2273_), .Y(_2274_) );
	OAI22X1 OAI22X1_186 ( .A(_2161_), .B(_2471__bF_buf13), .C(_2473__bF_buf7), .D(_2274_), .Y(_1002_) );
	OAI21X1 OAI21X1_585 ( .A(_1451_), .B(micro_hash_synth_W_9__1_), .C(_2231_), .Y(_2275_) );
	AOI21X1 AOI21X1_391 ( .A(micro_hash_synth_W_9__1_), .B(_1451_), .C(_2275_), .Y(_2276_) );
	OAI22X1 OAI22X1_187 ( .A(_1473_), .B(_2471__bF_buf12), .C(_2473__bF_buf6), .D(_2276_), .Y(_1004_) );
	OAI21X1 OAI21X1_586 ( .A(_1560_), .B(micro_hash_synth_W_9__2_), .C(_2233_), .Y(_2277_) );
	AOI21X1 AOI21X1_392 ( .A(micro_hash_synth_W_9__2_), .B(_1560_), .C(_2277_), .Y(_2278_) );
	OAI22X1 OAI22X1_188 ( .A(_2168_), .B(_2471__bF_buf11), .C(_2473__bF_buf5), .D(_2278_), .Y(_1005_) );
	OAI21X1 OAI21X1_587 ( .A(_1632_), .B(micro_hash_synth_W_9__3_), .C(_2235_), .Y(_2279_) );
	AOI21X1 AOI21X1_393 ( .A(micro_hash_synth_W_9__3_), .B(_1632_), .C(_2279_), .Y(_2280_) );
	OAI22X1 OAI22X1_189 ( .A(_1607_), .B(_2471__bF_buf10), .C(_2473__bF_buf4), .D(_2280_), .Y(_1006_) );
	OAI21X1 OAI21X1_588 ( .A(_1729_), .B(micro_hash_synth_W_9__4_), .C(_2237_), .Y(_2281_) );
	AOI21X1 AOI21X1_394 ( .A(micro_hash_synth_W_9__4_), .B(_1729_), .C(_2281_), .Y(_2282_) );
	OAI22X1 OAI22X1_190 ( .A(_1700_), .B(_2471__bF_buf9), .C(_2473__bF_buf3), .D(_2282_), .Y(_1007_) );
	OAI21X1 OAI21X1_589 ( .A(_2044_), .B(micro_hash_synth_W_9__5_), .C(_2239_), .Y(_2283_) );
	AOI21X1 AOI21X1_395 ( .A(micro_hash_synth_W_9__5_), .B(_2044_), .C(_2283_), .Y(_2284_) );
	OAI22X1 OAI22X1_191 ( .A(_2178_), .B(_2471__bF_buf8), .C(_2473__bF_buf2), .D(_2284_), .Y(_1008_) );
	OAI21X1 OAI21X1_590 ( .A(_2046_), .B(micro_hash_synth_W_9__6_), .C(_2241_), .Y(_2285_) );
	AOI21X1 AOI21X1_396 ( .A(micro_hash_synth_W_9__6_), .B(_2046_), .C(_2285_), .Y(_2286_) );
	OAI22X1 OAI22X1_192 ( .A(_2182_), .B(_2471__bF_buf7), .C(_2473__bF_buf1), .D(_2286_), .Y(_1009_) );
	OAI21X1 OAI21X1_591 ( .A(_2048_), .B(micro_hash_synth_W_9__7_), .C(_2243_), .Y(_2287_) );
	AOI21X1 AOI21X1_397 ( .A(micro_hash_synth_W_9__7_), .B(_2048_), .C(_2287_), .Y(_2288_) );
	OAI22X1 OAI22X1_193 ( .A(_2186_), .B(_2471__bF_buf6), .C(_2473__bF_buf0), .D(_2288_), .Y(_1010_) );
	INVX1 INVX1_600 ( .A(bloque_in_96_), .Y(_2289_) );
	OAI22X1 OAI22X1_194 ( .A(_2530_), .B(_2471__bF_buf5), .C(_2473__bF_buf15), .D(_2289_), .Y(_1011_) );
	INVX1 INVX1_601 ( .A(bloque_in_97_), .Y(_2290_) );
	OAI22X1 OAI22X1_195 ( .A(_2535_), .B(_2471__bF_buf4), .C(_2473__bF_buf14), .D(_2290_), .Y(_1012_) );
	INVX1 INVX1_602 ( .A(bloque_in_98_), .Y(_2291_) );
	OAI22X1 OAI22X1_196 ( .A(_2540_), .B(_2471__bF_buf3), .C(_2473__bF_buf13), .D(_2291_), .Y(_1013_) );
	INVX1 INVX1_603 ( .A(bloque_in_99_), .Y(_2292_) );
	OAI22X1 OAI22X1_197 ( .A(_2545_), .B(_2471__bF_buf2), .C(_2473__bF_buf12), .D(_2292_), .Y(_1014_) );
	INVX1 INVX1_604 ( .A(bloque_in_100_), .Y(_2293_) );
	OAI22X1 OAI22X1_198 ( .A(_2550_), .B(_2471__bF_buf1), .C(_2473__bF_buf11), .D(_2293_), .Y(_1015_) );
	INVX1 INVX1_605 ( .A(bloque_in_101_), .Y(_2294_) );
	OAI22X1 OAI22X1_199 ( .A(_2555_), .B(_2471__bF_buf0), .C(_2473__bF_buf10), .D(_2294_), .Y(_1016_) );
	INVX1 INVX1_606 ( .A(bloque_in_102_), .Y(_2295_) );
	OAI22X1 OAI22X1_200 ( .A(_2560_), .B(_2471__bF_buf13), .C(_2473__bF_buf9), .D(_2295_), .Y(_1017_) );
	INVX1 INVX1_607 ( .A(bloque_in_103_), .Y(_2296_) );
	OAI22X1 OAI22X1_201 ( .A(_2565_), .B(_2471__bF_buf12), .C(_2473__bF_buf8), .D(_2296_), .Y(_1018_) );
	INVX1 INVX1_608 ( .A(bloque_in_56_), .Y(_2297_) );
	OAI22X1 OAI22X1_202 ( .A(_2160_), .B(_2471__bF_buf11), .C(_2473__bF_buf7), .D(_2297_), .Y(_1020_) );
	INVX1 INVX1_609 ( .A(bloque_in_57_), .Y(_2298_) );
	OAI22X1 OAI22X1_203 ( .A(_2164_), .B(_2471__bF_buf10), .C(_2473__bF_buf6), .D(_2298_), .Y(_1021_) );
	INVX1 INVX1_610 ( .A(bloque_in_58_), .Y(_2299_) );
	OAI22X1 OAI22X1_204 ( .A(_2167_), .B(_2471__bF_buf9), .C(_2473__bF_buf5), .D(_2299_), .Y(_1022_) );
	INVX1 INVX1_611 ( .A(bloque_in_59_), .Y(_2300_) );
	OAI22X1 OAI22X1_205 ( .A(_2171_), .B(_2471__bF_buf8), .C(_2473__bF_buf4), .D(_2300_), .Y(_1023_) );
	INVX1 INVX1_612 ( .A(bloque_in_60_), .Y(_2301_) );
	OAI22X1 OAI22X1_206 ( .A(_2174_), .B(_2471__bF_buf7), .C(_2473__bF_buf3), .D(_2301_), .Y(_1024_) );
	INVX1 INVX1_613 ( .A(bloque_in_61_), .Y(_2302_) );
	OAI22X1 OAI22X1_207 ( .A(_2177_), .B(_2471__bF_buf6), .C(_2473__bF_buf2), .D(_2302_), .Y(_1025_) );
	INVX1 INVX1_614 ( .A(bloque_in_62_), .Y(_2303_) );
	OAI22X1 OAI22X1_208 ( .A(_2181_), .B(_2471__bF_buf5), .C(_2473__bF_buf1), .D(_2303_), .Y(_1026_) );
	INVX1 INVX1_615 ( .A(bloque_in_63_), .Y(_2304_) );
	OAI22X1 OAI22X1_209 ( .A(_2185_), .B(_2471__bF_buf4), .C(_2473__bF_buf0), .D(_2304_), .Y(_1027_) );
	INVX1 INVX1_616 ( .A(micro_hash_synth_W_14__0_), .Y(_2305_) );
	INVX1 INVX1_617 ( .A(bloque_in_112_), .Y(_2306_) );
	OAI22X1 OAI22X1_210 ( .A(_2305_), .B(_2471__bF_buf3), .C(_2473__bF_buf15), .D(_2306_), .Y(_1028_) );
	INVX1 INVX1_618 ( .A(bloque_in_113_), .Y(_2307_) );
	OAI22X1 OAI22X1_211 ( .A(_1501_), .B(_2471__bF_buf2), .C(_2473__bF_buf14), .D(_2307_), .Y(_1029_) );
	INVX1 INVX1_619 ( .A(micro_hash_synth_W_14__2_), .Y(_2308_) );
	INVX1 INVX1_620 ( .A(bloque_in_114_), .Y(_2309_) );
	OAI22X1 OAI22X1_212 ( .A(_2308_), .B(_2471__bF_buf1), .C(_2473__bF_buf13), .D(_2309_), .Y(_1030_) );
	INVX1 INVX1_621 ( .A(bloque_in_115_), .Y(_2310_) );
	OAI22X1 OAI22X1_213 ( .A(_1644_), .B(_2471__bF_buf0), .C(_2473__bF_buf12), .D(_2310_), .Y(_1031_) );
	INVX1 INVX1_622 ( .A(bloque_in_116_), .Y(_2311_) );
	OAI22X1 OAI22X1_214 ( .A(_1741_), .B(_2471__bF_buf13), .C(_2473__bF_buf11), .D(_2311_), .Y(_1032_) );
	INVX1 INVX1_623 ( .A(micro_hash_synth_W_14__5_), .Y(_2312_) );
	INVX1 INVX1_624 ( .A(bloque_in_117_), .Y(_2313_) );
	OAI22X1 OAI22X1_215 ( .A(_2312_), .B(_2471__bF_buf12), .C(_2473__bF_buf10), .D(_2313_), .Y(_1033_) );
	INVX1 INVX1_625 ( .A(micro_hash_synth_W_14__6_), .Y(_2314_) );
	INVX1 INVX1_626 ( .A(bloque_in_118_), .Y(_2315_) );
	OAI22X1 OAI22X1_216 ( .A(_2314_), .B(_2471__bF_buf11), .C(_2473__bF_buf9), .D(_2315_), .Y(_1034_) );
	INVX1 INVX1_627 ( .A(micro_hash_synth_W_14__7_), .Y(_2316_) );
	INVX1 INVX1_628 ( .A(bloque_in_119_), .Y(_2317_) );
	OAI22X1 OAI22X1_217 ( .A(_2316_), .B(_2471__bF_buf10), .C(_2473__bF_buf8), .D(_2317_), .Y(_1036_) );
	OAI21X1 OAI21X1_592 ( .A(_2030_), .B(micro_hash_synth_W_8__0_), .C(_2305_), .Y(_2318_) );
	AOI21X1 AOI21X1_398 ( .A(_2030_), .B(micro_hash_synth_W_8__0_), .C(_2318_), .Y(_2319_) );
	OAI22X1 OAI22X1_218 ( .A(_2196_), .B(_2471__bF_buf9), .C(_2473__bF_buf7), .D(_2319_), .Y(_1037_) );
	OAI21X1 OAI21X1_593 ( .A(_2031_), .B(micro_hash_synth_W_8__1_), .C(_1501_), .Y(_2320_) );
	AOI21X1 AOI21X1_399 ( .A(_2031_), .B(micro_hash_synth_W_8__1_), .C(_2320_), .Y(_2321_) );
	OAI22X1 OAI22X1_219 ( .A(_1432_), .B(_2471__bF_buf8), .C(_2473__bF_buf6), .D(_2321_), .Y(_1038_) );
	OAI21X1 OAI21X1_594 ( .A(_2032_), .B(micro_hash_synth_W_8__2_), .C(_2308_), .Y(_2322_) );
	AOI21X1 AOI21X1_400 ( .A(_2032_), .B(micro_hash_synth_W_8__2_), .C(_2322_), .Y(_2323_) );
	OAI22X1 OAI22X1_220 ( .A(_1529_), .B(_2471__bF_buf7), .C(_2473__bF_buf5), .D(_2323_), .Y(_1039_) );
	OAI21X1 OAI21X1_595 ( .A(_2033_), .B(micro_hash_synth_W_8__3_), .C(_1644_), .Y(_2324_) );
	AOI21X1 AOI21X1_401 ( .A(_2033_), .B(micro_hash_synth_W_8__3_), .C(_2324_), .Y(_2325_) );
	OAI22X1 OAI22X1_221 ( .A(_2203_), .B(_2471__bF_buf6), .C(_2473__bF_buf4), .D(_2325_), .Y(_1040_) );
	OAI21X1 OAI21X1_596 ( .A(_2034_), .B(micro_hash_synth_W_8__4_), .C(_1741_), .Y(_2326_) );
	AOI21X1 AOI21X1_402 ( .A(_2034_), .B(micro_hash_synth_W_8__4_), .C(_2326_), .Y(_2327_) );
	OAI22X1 OAI22X1_222 ( .A(_2206_), .B(_2471__bF_buf5), .C(_2473__bF_buf3), .D(_2327_), .Y(_1041_) );
	OAI21X1 OAI21X1_597 ( .A(_2035_), .B(micro_hash_synth_W_8__5_), .C(_2312_), .Y(_2328_) );
	AOI21X1 AOI21X1_403 ( .A(_2035_), .B(micro_hash_synth_W_8__5_), .C(_2328_), .Y(_2329_) );
	OAI22X1 OAI22X1_223 ( .A(_2210_), .B(_2471__bF_buf4), .C(_2473__bF_buf2), .D(_2329_), .Y(_1042_) );
	OAI21X1 OAI21X1_598 ( .A(_2036_), .B(micro_hash_synth_W_8__6_), .C(_2314_), .Y(_2330_) );
	AOI21X1 AOI21X1_404 ( .A(_2036_), .B(micro_hash_synth_W_8__6_), .C(_2330_), .Y(_2331_) );
	OAI22X1 OAI22X1_224 ( .A(_2214_), .B(_2471__bF_buf3), .C(_2473__bF_buf1), .D(_2331_), .Y(_1043_) );
	OAI21X1 OAI21X1_599 ( .A(_2037_), .B(micro_hash_synth_W_8__7_), .C(_2316_), .Y(_2332_) );
	AOI21X1 AOI21X1_405 ( .A(_2037_), .B(micro_hash_synth_W_8__7_), .C(_2332_), .Y(_2333_) );
	OAI22X1 OAI22X1_225 ( .A(_2218_), .B(_2471__bF_buf2), .C(_2473__bF_buf0), .D(_2333_), .Y(_1044_) );
	INVX1 INVX1_629 ( .A(micro_hash_synth_W_2__0_), .Y(_2334_) );
	OAI22X1 OAI22X1_226 ( .A(_2334_), .B(_2471__bF_buf1), .C(_2473__bF_buf15), .D(_1956_), .Y(_1045_) );
	OAI22X1 OAI22X1_227 ( .A(_1496_), .B(_2471__bF_buf0), .C(_2473__bF_buf14), .D(_1957_), .Y(_1046_) );
	INVX1 INVX1_630 ( .A(micro_hash_synth_W_2__2_), .Y(_2335_) );
	OAI22X1 OAI22X1_228 ( .A(_2335_), .B(_2471__bF_buf13), .C(_2473__bF_buf13), .D(_1958_), .Y(_1047_) );
	OAI22X1 OAI22X1_229 ( .A(_1636_), .B(_2471__bF_buf12), .C(_2473__bF_buf12), .D(_1959_), .Y(_1048_) );
	OAI22X1 OAI22X1_230 ( .A(_1733_), .B(_2471__bF_buf11), .C(_2473__bF_buf11), .D(_1960_), .Y(_1049_) );
	INVX1 INVX1_631 ( .A(micro_hash_synth_W_2__5_), .Y(_2336_) );
	OAI22X1 OAI22X1_231 ( .A(_2336_), .B(_2471__bF_buf10), .C(_2473__bF_buf10), .D(_1961_), .Y(_1050_) );
	INVX1 INVX1_632 ( .A(micro_hash_synth_W_2__6_), .Y(_2337_) );
	OAI22X1 OAI22X1_232 ( .A(_2337_), .B(_2471__bF_buf9), .C(_2473__bF_buf9), .D(_1962_), .Y(_1051_) );
	INVX1 INVX1_633 ( .A(micro_hash_synth_W_2__7_), .Y(_2338_) );
	OAI22X1 OAI22X1_233 ( .A(_2338_), .B(_2471__bF_buf8), .C(_2473__bF_buf8), .D(_1963_), .Y(_1052_) );
	INVX1 INVX1_634 ( .A(bloque_in_104_), .Y(_2339_) );
	OAI22X1 OAI22X1_234 ( .A(_2474_), .B(_2471__bF_buf7), .C(_2473__bF_buf7), .D(_2339_), .Y(_1053_) );
	INVX1 INVX1_635 ( .A(bloque_in_105_), .Y(_2340_) );
	OAI22X1 OAI22X1_235 ( .A(_2479_), .B(_2471__bF_buf6), .C(_2473__bF_buf6), .D(_2340_), .Y(_1054_) );
	INVX1 INVX1_636 ( .A(bloque_in_106_), .Y(_2341_) );
	OAI22X1 OAI22X1_236 ( .A(_2484_), .B(_2471__bF_buf5), .C(_2473__bF_buf5), .D(_2341_), .Y(_1055_) );
	INVX1 INVX1_637 ( .A(bloque_in_107_), .Y(_2342_) );
	OAI22X1 OAI22X1_237 ( .A(_2489_), .B(_2471__bF_buf4), .C(_2473__bF_buf4), .D(_2342_), .Y(_1056_) );
	INVX1 INVX1_638 ( .A(bloque_in_108_), .Y(_2343_) );
	OAI22X1 OAI22X1_238 ( .A(_2494_), .B(_2471__bF_buf3), .C(_2473__bF_buf3), .D(_2343_), .Y(_1057_) );
	INVX1 INVX1_639 ( .A(bloque_in_109_), .Y(_2344_) );
	OAI22X1 OAI22X1_239 ( .A(_2499_), .B(_2471__bF_buf2), .C(_2473__bF_buf2), .D(_2344_), .Y(_1058_) );
	INVX1 INVX1_640 ( .A(bloque_in_110_), .Y(_2345_) );
	OAI22X1 OAI22X1_240 ( .A(_2504_), .B(_2471__bF_buf1), .C(_2473__bF_buf1), .D(_2345_), .Y(_1059_) );
	INVX1 INVX1_641 ( .A(bloque_in_111_), .Y(_2346_) );
	OAI22X1 OAI22X1_241 ( .A(_2509_), .B(_2471__bF_buf0), .C(_2473__bF_buf0), .D(_2346_), .Y(_1060_) );
	OAI21X1 OAI21X1_600 ( .A(_2334_), .B(micro_hash_synth_W_7__0_), .C(_2474_), .Y(_2347_) );
	AOI21X1 AOI21X1_406 ( .A(_2334_), .B(micro_hash_synth_W_7__0_), .C(_2347_), .Y(_2348_) );
	OAI22X1 OAI22X1_242 ( .A(_2245_), .B(_2471__bF_buf13), .C(_2473__bF_buf15), .D(_2348_), .Y(_1061_) );
	OAI21X1 OAI21X1_601 ( .A(_1496_), .B(micro_hash_synth_W_7__1_), .C(_2479_), .Y(_2349_) );
	AOI21X1 AOI21X1_407 ( .A(_1496_), .B(micro_hash_synth_W_7__1_), .C(_2349_), .Y(_2350_) );
	OAI22X1 OAI22X1_243 ( .A(_1429_), .B(_2471__bF_buf12), .C(_2473__bF_buf14), .D(_2350_), .Y(_1062_) );
	OAI21X1 OAI21X1_602 ( .A(_2335_), .B(micro_hash_synth_W_7__2_), .C(_2484_), .Y(_2351_) );
	AOI21X1 AOI21X1_408 ( .A(_2335_), .B(micro_hash_synth_W_7__2_), .C(_2351_), .Y(_2352_) );
	OAI22X1 OAI22X1_244 ( .A(_1527_), .B(_2471__bF_buf11), .C(_2473__bF_buf13), .D(_2352_), .Y(_1063_) );
	OAI21X1 OAI21X1_603 ( .A(_1636_), .B(micro_hash_synth_W_7__3_), .C(_2489_), .Y(_2353_) );
	AOI21X1 AOI21X1_409 ( .A(_1636_), .B(micro_hash_synth_W_7__3_), .C(_2353_), .Y(_2354_) );
	OAI22X1 OAI22X1_245 ( .A(_1610_), .B(_2471__bF_buf10), .C(_2473__bF_buf12), .D(_2354_), .Y(_1064_) );
	OAI21X1 OAI21X1_604 ( .A(_1733_), .B(micro_hash_synth_W_7__4_), .C(_2494_), .Y(_2355_) );
	AOI21X1 AOI21X1_410 ( .A(_1733_), .B(micro_hash_synth_W_7__4_), .C(_2355_), .Y(_2356_) );
	OAI22X1 OAI22X1_246 ( .A(_1697_), .B(_2471__bF_buf9), .C(_2473__bF_buf11), .D(_2356_), .Y(_1065_) );
	OAI21X1 OAI21X1_605 ( .A(_2336_), .B(micro_hash_synth_W_7__5_), .C(_2499_), .Y(_2357_) );
	AOI21X1 AOI21X1_411 ( .A(_2336_), .B(micro_hash_synth_W_7__5_), .C(_2357_), .Y(_2358_) );
	OAI22X1 OAI22X1_247 ( .A(_2256_), .B(_2471__bF_buf8), .C(_2473__bF_buf10), .D(_2358_), .Y(_1066_) );
	OAI21X1 OAI21X1_606 ( .A(_2337_), .B(micro_hash_synth_W_7__6_), .C(_2504_), .Y(_2359_) );
	AOI21X1 AOI21X1_412 ( .A(_2337_), .B(micro_hash_synth_W_7__6_), .C(_2359_), .Y(_2360_) );
	OAI22X1 OAI22X1_248 ( .A(_2259_), .B(_2471__bF_buf7), .C(_2473__bF_buf9), .D(_2360_), .Y(_1067_) );
	OAI21X1 OAI21X1_607 ( .A(_2338_), .B(micro_hash_synth_W_7__7_), .C(_2509_), .Y(_2361_) );
	AOI21X1 AOI21X1_413 ( .A(_2338_), .B(micro_hash_synth_W_7__7_), .C(_2361_), .Y(_2362_) );
	OAI22X1 OAI22X1_249 ( .A(_2262_), .B(_2471__bF_buf6), .C(_2473__bF_buf8), .D(_2362_), .Y(_1068_) );
	INVX1 INVX1_642 ( .A(bloque_in_80_), .Y(_2363_) );
	OAI22X1 OAI22X1_250 ( .A(_2058_), .B(_2471__bF_buf5), .C(_2473__bF_buf7), .D(_2363_), .Y(_1069_) );
	INVX1 INVX1_643 ( .A(bloque_in_81_), .Y(_2364_) );
	OAI22X1 OAI22X1_251 ( .A(_1507_), .B(_2471__bF_buf4), .C(_2473__bF_buf6), .D(_2364_), .Y(_1070_) );
	INVX1 INVX1_644 ( .A(bloque_in_82_), .Y(_2365_) );
	OAI22X1 OAI22X1_252 ( .A(_2065_), .B(_2471__bF_buf3), .C(_2473__bF_buf5), .D(_2365_), .Y(_1071_) );
	INVX1 INVX1_645 ( .A(bloque_in_83_), .Y(_2366_) );
	OAI22X1 OAI22X1_253 ( .A(_1650_), .B(_2471__bF_buf2), .C(_2473__bF_buf4), .D(_2366_), .Y(_1072_) );
	INVX1 INVX1_646 ( .A(bloque_in_84_), .Y(_2367_) );
	OAI22X1 OAI22X1_254 ( .A(_1747_), .B(_2471__bF_buf1), .C(_2473__bF_buf3), .D(_2367_), .Y(_1073_) );
	INVX1 INVX1_647 ( .A(bloque_in_85_), .Y(_2368_) );
	OAI22X1 OAI22X1_255 ( .A(_2075_), .B(_2471__bF_buf0), .C(_2473__bF_buf2), .D(_2368_), .Y(_1074_) );
	INVX1 INVX1_648 ( .A(bloque_in_86_), .Y(_2369_) );
	OAI22X1 OAI22X1_256 ( .A(_2079_), .B(_2471__bF_buf13), .C(_2473__bF_buf1), .D(_2369_), .Y(_1075_) );
	INVX1 INVX1_649 ( .A(bloque_in_87_), .Y(_2370_) );
	OAI22X1 OAI22X1_257 ( .A(_2083_), .B(_2471__bF_buf12), .C(_2473__bF_buf0), .D(_2370_), .Y(_1076_) );
	INVX1 INVX1_650 ( .A(micro_hash_synth_W_28__0_), .Y(_2371_) );
	OAI21X1 OAI21X1_608 ( .A(_2305_), .B(micro_hash_synth_W_19__0_), .C(_2569_), .Y(_2372_) );
	AOI21X1 AOI21X1_414 ( .A(_2305_), .B(micro_hash_synth_W_19__0_), .C(_2372_), .Y(_2373_) );
	OAI22X1 OAI22X1_258 ( .A(_2371_), .B(_2471__bF_buf11), .C(_2473__bF_buf15), .D(_2373_), .Y(_1077_) );
	OAI21X1 OAI21X1_609 ( .A(_1501_), .B(micro_hash_synth_W_19__1_), .C(_2574_), .Y(_2374_) );
	AOI21X1 AOI21X1_415 ( .A(_1501_), .B(micro_hash_synth_W_19__1_), .C(_2374_), .Y(_2375_) );
	OAI22X1 OAI22X1_259 ( .A(_1438_), .B(_2471__bF_buf10), .C(_2473__bF_buf14), .D(_2375_), .Y(_1078_) );
	INVX1 INVX1_651 ( .A(micro_hash_synth_W_28__2_), .Y(_2376_) );
	OAI21X1 OAI21X1_610 ( .A(_2308_), .B(micro_hash_synth_W_19__2_), .C(_2579_), .Y(_2377_) );
	AOI21X1 AOI21X1_416 ( .A(_2308_), .B(micro_hash_synth_W_19__2_), .C(_2377_), .Y(_2378_) );
	OAI22X1 OAI22X1_260 ( .A(_2376_), .B(_2471__bF_buf9), .C(_2473__bF_buf13), .D(_2378_), .Y(_1079_) );
	OAI21X1 OAI21X1_611 ( .A(_1644_), .B(micro_hash_synth_W_19__3_), .C(_2584_), .Y(_2379_) );
	AOI21X1 AOI21X1_417 ( .A(_1644_), .B(micro_hash_synth_W_19__3_), .C(_2379_), .Y(_2380_) );
	OAI22X1 OAI22X1_261 ( .A(_1618_), .B(_2471__bF_buf8), .C(_2473__bF_buf12), .D(_2380_), .Y(_1080_) );
	OAI21X1 OAI21X1_612 ( .A(_1741_), .B(micro_hash_synth_W_19__4_), .C(_2589_), .Y(_2381_) );
	AOI21X1 AOI21X1_418 ( .A(_1741_), .B(micro_hash_synth_W_19__4_), .C(_2381_), .Y(_2382_) );
	OAI22X1 OAI22X1_262 ( .A(_1719_), .B(_2471__bF_buf7), .C(_2473__bF_buf11), .D(_2382_), .Y(_1081_) );
	INVX1 INVX1_652 ( .A(micro_hash_synth_W_28__5_), .Y(_2383_) );
	OAI21X1 OAI21X1_613 ( .A(_2312_), .B(micro_hash_synth_W_19__5_), .C(_2594_), .Y(_2384_) );
	AOI21X1 AOI21X1_419 ( .A(_2312_), .B(micro_hash_synth_W_19__5_), .C(_2384_), .Y(_2385_) );
	OAI22X1 OAI22X1_263 ( .A(_2383_), .B(_2471__bF_buf6), .C(_2473__bF_buf10), .D(_2385_), .Y(_1082_) );
	INVX1 INVX1_653 ( .A(micro_hash_synth_W_28__6_), .Y(_2386_) );
	OAI21X1 OAI21X1_614 ( .A(_2314_), .B(micro_hash_synth_W_19__6_), .C(_2599_), .Y(_2387_) );
	AOI21X1 AOI21X1_420 ( .A(_2314_), .B(micro_hash_synth_W_19__6_), .C(_2387_), .Y(_2388_) );
	OAI22X1 OAI22X1_264 ( .A(_2386_), .B(_2471__bF_buf5), .C(_2473__bF_buf9), .D(_2388_), .Y(_1083_) );
	INVX1 INVX1_654 ( .A(micro_hash_synth_W_28__7_), .Y(_2389_) );
	OAI21X1 OAI21X1_615 ( .A(_2316_), .B(micro_hash_synth_W_19__7_), .C(_2604_), .Y(_2390_) );
	AOI21X1 AOI21X1_421 ( .A(_2316_), .B(micro_hash_synth_W_19__7_), .C(_2390_), .Y(_2391_) );
	OAI22X1 OAI22X1_265 ( .A(_2389_), .B(_2471__bF_buf4), .C(_2473__bF_buf8), .D(_2391_), .Y(_1084_) );
	NAND2X1 NAND2X1_243 ( .A(micro_hash_synth_W_29__0_), .B(_2189__bF_buf1), .Y(_2392_) );
	OAI21X1 OAI21X1_616 ( .A(_2229_), .B(micro_hash_synth_W_20__0_), .C(_2529_), .Y(_2393_) );
	AOI21X1 AOI21X1_422 ( .A(_2229_), .B(micro_hash_synth_W_20__0_), .C(_2393_), .Y(_2394_) );
	OAI21X1 OAI21X1_617 ( .A(_2473__bF_buf7), .B(_2394_), .C(_2392_), .Y(_1085_) );
	NAND2X1 NAND2X1_244 ( .A(micro_hash_synth_W_29__1_), .B(_2189__bF_buf0), .Y(_2395_) );
	OAI21X1 OAI21X1_618 ( .A(_2231_), .B(micro_hash_synth_W_20__1_), .C(_2534_), .Y(_2396_) );
	AOI21X1 AOI21X1_423 ( .A(_2231_), .B(micro_hash_synth_W_20__1_), .C(_2396_), .Y(_2397_) );
	OAI21X1 OAI21X1_619 ( .A(_2473__bF_buf6), .B(_2397_), .C(_2395_), .Y(_1086_) );
	NAND2X1 NAND2X1_245 ( .A(micro_hash_synth_W_29__2_), .B(_2189__bF_buf4), .Y(_2398_) );
	OAI21X1 OAI21X1_620 ( .A(_2233_), .B(micro_hash_synth_W_20__2_), .C(_2539_), .Y(_2399_) );
	AOI21X1 AOI21X1_424 ( .A(_2233_), .B(micro_hash_synth_W_20__2_), .C(_2399_), .Y(_2400_) );
	OAI21X1 OAI21X1_621 ( .A(_2473__bF_buf5), .B(_2400_), .C(_2398_), .Y(_1087_) );
	NAND2X1 NAND2X1_246 ( .A(micro_hash_synth_W_29__3_), .B(_2189__bF_buf3), .Y(_2401_) );
	OAI21X1 OAI21X1_622 ( .A(_2235_), .B(micro_hash_synth_W_20__3_), .C(_2544_), .Y(_2402_) );
	AOI21X1 AOI21X1_425 ( .A(_2235_), .B(micro_hash_synth_W_20__3_), .C(_2402_), .Y(_2403_) );
	OAI21X1 OAI21X1_623 ( .A(_2473__bF_buf4), .B(_2403_), .C(_2401_), .Y(_1088_) );
	NAND2X1 NAND2X1_247 ( .A(micro_hash_synth_W_29__4_), .B(_2189__bF_buf2), .Y(_2404_) );
	OAI21X1 OAI21X1_624 ( .A(_2237_), .B(micro_hash_synth_W_20__4_), .C(_2549_), .Y(_2405_) );
	AOI21X1 AOI21X1_426 ( .A(_2237_), .B(micro_hash_synth_W_20__4_), .C(_2405_), .Y(_2406_) );
	OAI21X1 OAI21X1_625 ( .A(_2473__bF_buf3), .B(_2406_), .C(_2404_), .Y(_1089_) );
	NAND2X1 NAND2X1_248 ( .A(micro_hash_synth_W_29__5_), .B(_2189__bF_buf1), .Y(_2407_) );
	OAI21X1 OAI21X1_626 ( .A(_2239_), .B(micro_hash_synth_W_20__5_), .C(_2554_), .Y(_2408_) );
	AOI21X1 AOI21X1_427 ( .A(_2239_), .B(micro_hash_synth_W_20__5_), .C(_2408_), .Y(_2409_) );
	OAI21X1 OAI21X1_627 ( .A(_2473__bF_buf2), .B(_2409_), .C(_2407_), .Y(_1090_) );
	NAND2X1 NAND2X1_249 ( .A(micro_hash_synth_W_29__6_), .B(_2189__bF_buf0), .Y(_2410_) );
	OAI21X1 OAI21X1_628 ( .A(_2241_), .B(micro_hash_synth_W_20__6_), .C(_2559_), .Y(_2411_) );
	AOI21X1 AOI21X1_428 ( .A(_2241_), .B(micro_hash_synth_W_20__6_), .C(_2411_), .Y(_2412_) );
	OAI21X1 OAI21X1_629 ( .A(_2473__bF_buf1), .B(_2412_), .C(_2410_), .Y(_1091_) );
	NAND2X1 NAND2X1_250 ( .A(micro_hash_synth_W_29__7_), .B(_2189__bF_buf4), .Y(_2413_) );
	OAI21X1 OAI21X1_630 ( .A(_2243_), .B(micro_hash_synth_W_20__7_), .C(_2564_), .Y(_2414_) );
	AOI21X1 AOI21X1_429 ( .A(_2243_), .B(micro_hash_synth_W_20__7_), .C(_2414_), .Y(_2415_) );
	OAI21X1 OAI21X1_631 ( .A(_2473__bF_buf0), .B(_2415_), .C(_2413_), .Y(_1092_) );
	NAND2X1 NAND2X1_251 ( .A(micro_hash_synth_W_30__0_), .B(_2189__bF_buf3), .Y(_2416_) );
	OAI21X1 OAI21X1_632 ( .A(_2245_), .B(micro_hash_synth_W_21__0_), .C(_2461_), .Y(_2417_) );
	AOI21X1 AOI21X1_430 ( .A(_2245_), .B(micro_hash_synth_W_21__0_), .C(_2417_), .Y(_2418_) );
	OAI21X1 OAI21X1_633 ( .A(_2473__bF_buf15), .B(_2418_), .C(_2416_), .Y(_1093_) );
	OAI21X1 OAI21X1_634 ( .A(_1429_), .B(micro_hash_synth_W_21__1_), .C(_2478_), .Y(_2419_) );
	AOI21X1 AOI21X1_431 ( .A(_1429_), .B(micro_hash_synth_W_21__1_), .C(_2419_), .Y(_2420_) );
	OAI22X1 OAI22X1_266 ( .A(_1441_), .B(_2471__bF_buf3), .C(_2473__bF_buf14), .D(_2420_), .Y(_1094_) );
	NAND2X1 NAND2X1_252 ( .A(micro_hash_synth_W_30__2_), .B(_2189__bF_buf2), .Y(_2421_) );
	OAI21X1 OAI21X1_635 ( .A(_1527_), .B(micro_hash_synth_W_21__2_), .C(_2483_), .Y(_2422_) );
	AOI21X1 AOI21X1_432 ( .A(_1527_), .B(micro_hash_synth_W_21__2_), .C(_2422_), .Y(_2423_) );
	OAI21X1 OAI21X1_636 ( .A(_2473__bF_buf13), .B(_2423_), .C(_2421_), .Y(_1095_) );
	OAI21X1 OAI21X1_637 ( .A(_1610_), .B(micro_hash_synth_W_21__3_), .C(_2488_), .Y(_2424_) );
	AOI21X1 AOI21X1_433 ( .A(_1610_), .B(micro_hash_synth_W_21__3_), .C(_2424_), .Y(_2425_) );
	OAI22X1 OAI22X1_267 ( .A(_1615_), .B(_2471__bF_buf2), .C(_2473__bF_buf12), .D(_2425_), .Y(_1096_) );
	OAI21X1 OAI21X1_638 ( .A(_1697_), .B(micro_hash_synth_W_21__4_), .C(_2493_), .Y(_2426_) );
	AOI21X1 AOI21X1_434 ( .A(_1697_), .B(micro_hash_synth_W_21__4_), .C(_2426_), .Y(_2427_) );
	OAI22X1 OAI22X1_268 ( .A(_1716_), .B(_2471__bF_buf1), .C(_2473__bF_buf11), .D(_2427_), .Y(_1097_) );
	NAND2X1 NAND2X1_253 ( .A(micro_hash_synth_W_30__5_), .B(_2189__bF_buf1), .Y(_2428_) );
	OAI21X1 OAI21X1_639 ( .A(_2256_), .B(micro_hash_synth_W_21__5_), .C(_2498_), .Y(_2429_) );
	AOI21X1 AOI21X1_435 ( .A(_2256_), .B(micro_hash_synth_W_21__5_), .C(_2429_), .Y(_2430_) );
	OAI21X1 OAI21X1_640 ( .A(_2473__bF_buf10), .B(_2430_), .C(_2428_), .Y(_1098_) );
	NAND2X1 NAND2X1_254 ( .A(micro_hash_synth_W_30__6_), .B(_2189__bF_buf0), .Y(_2431_) );
	OAI21X1 OAI21X1_641 ( .A(_2259_), .B(micro_hash_synth_W_21__6_), .C(_2503_), .Y(_2432_) );
	AOI21X1 AOI21X1_436 ( .A(_2259_), .B(micro_hash_synth_W_21__6_), .C(_2432_), .Y(_2433_) );
	OAI21X1 OAI21X1_642 ( .A(_2473__bF_buf9), .B(_2433_), .C(_2431_), .Y(_1099_) );
	NAND2X1 NAND2X1_255 ( .A(micro_hash_synth_W_30__7_), .B(_2189__bF_buf4), .Y(_2434_) );
	OAI21X1 OAI21X1_643 ( .A(_2262_), .B(micro_hash_synth_W_21__7_), .C(_2508_), .Y(_2435_) );
	AOI21X1 AOI21X1_437 ( .A(_2262_), .B(micro_hash_synth_W_21__7_), .C(_2435_), .Y(_2436_) );
	OAI21X1 OAI21X1_644 ( .A(_2473__bF_buf8), .B(_2436_), .C(_2434_), .Y(_1100_) );
	NAND2X1 NAND2X1_256 ( .A(micro_hash_synth_W_31__0_), .B(_2189__bF_buf3), .Y(_2437_) );
	OAI21X1 OAI21X1_645 ( .A(_2196_), .B(micro_hash_synth_W_22__0_), .C(_2371_), .Y(_2438_) );
	AOI21X1 AOI21X1_438 ( .A(_2196_), .B(micro_hash_synth_W_22__0_), .C(_2438_), .Y(_2439_) );
	OAI21X1 OAI21X1_646 ( .A(_2473__bF_buf7), .B(_2439_), .C(_2437_), .Y(_1101_) );
	NAND2X1 NAND2X1_257 ( .A(micro_hash_synth_W_31__1_), .B(_2189__bF_buf2), .Y(_2440_) );
	OAI21X1 OAI21X1_647 ( .A(_1432_), .B(micro_hash_synth_W_22__1_), .C(_1438_), .Y(_2441_) );
	AOI21X1 AOI21X1_439 ( .A(_1432_), .B(micro_hash_synth_W_22__1_), .C(_2441_), .Y(_2442_) );
	OAI21X1 OAI21X1_648 ( .A(_2473__bF_buf6), .B(_2442_), .C(_2440_), .Y(_1102_) );
	NAND2X1 NAND2X1_258 ( .A(micro_hash_synth_W_31__2_), .B(_2189__bF_buf1), .Y(_2443_) );
	OAI21X1 OAI21X1_649 ( .A(_1529_), .B(micro_hash_synth_W_22__2_), .C(_2376_), .Y(_2444_) );
	AOI21X1 AOI21X1_440 ( .A(_1529_), .B(micro_hash_synth_W_22__2_), .C(_2444_), .Y(_2445_) );
	OAI21X1 OAI21X1_650 ( .A(_2473__bF_buf5), .B(_2445_), .C(_2443_), .Y(_1103_) );
	NAND2X1 NAND2X1_259 ( .A(micro_hash_synth_W_31__3_), .B(_2189__bF_buf0), .Y(_2446_) );
	OAI21X1 OAI21X1_651 ( .A(_2203_), .B(micro_hash_synth_W_22__3_), .C(_1618_), .Y(_2447_) );
	AOI21X1 AOI21X1_441 ( .A(_2203_), .B(micro_hash_synth_W_22__3_), .C(_2447_), .Y(_2448_) );
	OAI21X1 OAI21X1_652 ( .A(_2473__bF_buf4), .B(_2448_), .C(_2446_), .Y(_1104_) );
	NAND2X1 NAND2X1_260 ( .A(micro_hash_synth_W_31__4_), .B(_2189__bF_buf4), .Y(_2449_) );
	OAI21X1 OAI21X1_653 ( .A(_2206_), .B(micro_hash_synth_W_22__4_), .C(_1719_), .Y(_2450_) );
	AOI21X1 AOI21X1_442 ( .A(_2206_), .B(micro_hash_synth_W_22__4_), .C(_2450_), .Y(_2451_) );
	OAI21X1 OAI21X1_654 ( .A(_2473__bF_buf3), .B(_2451_), .C(_2449_), .Y(_1105_) );
	NAND2X1 NAND2X1_261 ( .A(micro_hash_synth_W_31__5_), .B(_2189__bF_buf3), .Y(_2452_) );
	OAI21X1 OAI21X1_655 ( .A(_2210_), .B(micro_hash_synth_W_22__5_), .C(_2383_), .Y(_2453_) );
	AOI21X1 AOI21X1_443 ( .A(_2210_), .B(micro_hash_synth_W_22__5_), .C(_2453_), .Y(_2454_) );
	OAI21X1 OAI21X1_656 ( .A(_2473__bF_buf2), .B(_2454_), .C(_2452_), .Y(_1106_) );
	NAND2X1 NAND2X1_262 ( .A(micro_hash_synth_W_31__6_), .B(_2189__bF_buf2), .Y(_2455_) );
	OAI21X1 OAI21X1_657 ( .A(_2214_), .B(micro_hash_synth_W_22__6_), .C(_2386_), .Y(_2456_) );
	AOI21X1 AOI21X1_444 ( .A(_2214_), .B(micro_hash_synth_W_22__6_), .C(_2456_), .Y(_2457_) );
	OAI21X1 OAI21X1_658 ( .A(_2473__bF_buf1), .B(_2457_), .C(_2455_), .Y(_1107_) );
	NAND2X1 NAND2X1_263 ( .A(micro_hash_synth_W_31__7_), .B(_2189__bF_buf1), .Y(_2458_) );
	OAI21X1 OAI21X1_659 ( .A(_2218_), .B(micro_hash_synth_W_22__7_), .C(_2389_), .Y(_2459_) );
	AOI21X1 AOI21X1_445 ( .A(_2218_), .B(micro_hash_synth_W_22__7_), .C(_2459_), .Y(_2460_) );
	OAI21X1 OAI21X1_660 ( .A(_2473__bF_buf0), .B(_2460_), .C(_2458_), .Y(_1108_) );
	DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf44), .D(_1167_), .Q(micro_hash_synth_W_22__0_) );
	DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf43), .D(_1168_), .Q(micro_hash_synth_W_22__1_) );
	DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf42), .D(_1170_), .Q(micro_hash_synth_W_22__2_) );
	DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf41), .D(_1171_), .Q(micro_hash_synth_W_22__3_) );
	DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf40), .D(_1172_), .Q(micro_hash_synth_W_22__4_) );
	DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf39), .D(_1173_), .Q(micro_hash_synth_W_22__5_) );
	DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf38), .D(_1174_), .Q(micro_hash_synth_W_22__6_) );
	DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf37), .D(_1175_), .Q(micro_hash_synth_W_22__7_) );
	DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf36), .D(_951_), .Q(micro_hash_synth_W_0__0_) );
	DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf35), .D(_952_), .Q(micro_hash_synth_W_0__1_) );
	DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf34), .D(_953_), .Q(micro_hash_synth_W_0__2_) );
	DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf33), .D(_954_), .Q(micro_hash_synth_W_0__3_) );
	DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf32), .D(_956_), .Q(micro_hash_synth_W_0__4_) );
	DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf31), .D(_957_), .Q(micro_hash_synth_W_0__5_) );
	DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf30), .D(_958_), .Q(micro_hash_synth_W_0__6_) );
	DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf29), .D(_959_), .Q(micro_hash_synth_W_0__7_) );
	DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf28), .D(_942_), .Q(micro_hash_synth_W_21__0_) );
	DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf27), .D(_943_), .Q(micro_hash_synth_W_21__1_) );
	DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf26), .D(_944_), .Q(micro_hash_synth_W_21__2_) );
	DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf25), .D(_945_), .Q(micro_hash_synth_W_21__3_) );
	DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf24), .D(_946_), .Q(micro_hash_synth_W_21__4_) );
	DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf23), .D(_947_), .Q(micro_hash_synth_W_21__5_) );
	DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf22), .D(_948_), .Q(micro_hash_synth_W_21__6_) );
	DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf21), .D(_949_), .Q(micro_hash_synth_W_21__7_) );
	DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf20), .D(_960_), .Q(micro_hash_synth_W_20__0_) );
	DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf19), .D(_961_), .Q(micro_hash_synth_W_20__1_) );
	DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf18), .D(_962_), .Q(micro_hash_synth_W_20__2_) );
	DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_bF_buf17), .D(_963_), .Q(micro_hash_synth_W_20__3_) );
	DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_bF_buf16), .D(_964_), .Q(micro_hash_synth_W_20__4_) );
	DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_bF_buf15), .D(_965_), .Q(micro_hash_synth_W_20__5_) );
	DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_bF_buf14), .D(_966_), .Q(micro_hash_synth_W_20__6_) );
	DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_bF_buf13), .D(_967_), .Q(micro_hash_synth_W_20__7_) );
	DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_bF_buf12), .D(_985_), .Q(micro_hash_synth_W_19__0_) );
	DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_bF_buf11), .D(_986_), .Q(micro_hash_synth_W_19__1_) );
	DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_bF_buf10), .D(_988_), .Q(micro_hash_synth_W_19__2_) );
	DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_bF_buf9), .D(_989_), .Q(micro_hash_synth_W_19__3_) );
	DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_bF_buf8), .D(_990_), .Q(micro_hash_synth_W_19__4_) );
	DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_bF_buf7), .D(_991_), .Q(micro_hash_synth_W_19__5_) );
	DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_bF_buf6), .D(_992_), .Q(micro_hash_synth_W_19__6_) );
	DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_bF_buf5), .D(_993_), .Q(micro_hash_synth_W_19__7_) );
	DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_bF_buf4), .D(_927__0_), .Q(H_0_) );
	DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_bF_buf3), .D(_927__1_), .Q(H_1_) );
	DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_bF_buf2), .D(_927__2_), .Q(H_2_) );
	DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_bF_buf1), .D(_927__3_), .Q(H_3_) );
	DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_bF_buf0), .D(_927__4_), .Q(H_4_) );
	DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_bF_buf76), .D(_927__5_), .Q(H_5_) );
	DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_bF_buf75), .D(_927__6_), .Q(H_6_) );
	DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_bF_buf74), .D(_927__7_), .Q(H_7_) );
	DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_bF_buf73), .D(_927__8_), .Q(H_8_) );
	DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_bF_buf72), .D(_927__9_), .Q(H_9_) );
	DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_bF_buf71), .D(_927__10_), .Q(H_10_) );
	DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_bF_buf70), .D(_927__11_), .Q(H_11_) );
	DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_bF_buf69), .D(_927__12_), .Q(H_12_) );
	DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_bF_buf68), .D(_927__13_), .Q(H_13_) );
	DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_bF_buf67), .D(_927__14_), .Q(H_14_) );
	DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_bF_buf66), .D(_927__15_), .Q(H_15_) );
	DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_bF_buf65), .D(_927__16_), .Q(H_16_) );
	DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_bF_buf64), .D(_927__17_), .Q(H_17_) );
	DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_bF_buf63), .D(_927__18_), .Q(H_18_) );
	DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_bF_buf62), .D(_927__19_), .Q(H_19_) );
	DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_bF_buf61), .D(_927__20_), .Q(H_20_) );
	DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_bF_buf60), .D(_927__21_), .Q(H_21_) );
	DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_bF_buf59), .D(_927__22_), .Q(H_22_) );
	DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_bF_buf58), .D(_927__23_), .Q(H_23_) );
	DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_bF_buf57), .D(_931__0_), .Q(concatenador_count_0_) );
	DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_bF_buf56), .D(_931__1_), .Q(concatenador_count_1_) );
	DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_bF_buf55), .D(_931__2_), .Q(concatenador_count_2_) );
	DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_bF_buf54), .D(_931__3_), .Q(concatenador_count_3_) );
	DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_bF_buf53), .D(_931__4_), .Q(concatenador_count_4_) );
	DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_bF_buf52), .D(_931__5_), .Q(concatenador_count_5_) );
	DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_bF_buf51), .D(_933__0_), .Q(comparador_nonce_synth_1_0_) );
	DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_bF_buf50), .D(_933__1_), .Q(comparador_nonce_synth_1_1_) );
	DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_bF_buf49), .D(_933__2_), .Q(comparador_nonce_synth_1_2_) );
	DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_bF_buf48), .D(_933__3_), .Q(comparador_nonce_synth_1_3_) );
	DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_bF_buf47), .D(_933__4_), .Q(comparador_nonce_synth_1_4_) );
	DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_bF_buf46), .D(_933__5_), .Q(comparador_nonce_synth_1_5_) );
	DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_bF_buf45), .D(_933__6_), .Q(comparador_nonce_synth_1_6_) );
	DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_bF_buf44), .D(_933__7_), .Q(comparador_nonce_synth_1_7_) );
	DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_bF_buf43), .D(_933__8_), .Q(comparador_nonce_synth_1_8_) );
	DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_bF_buf42), .D(_933__9_), .Q(comparador_nonce_synth_1_9_) );
	DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_bF_buf41), .D(_933__10_), .Q(comparador_nonce_synth_1_10_) );
	DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_bF_buf40), .D(_933__11_), .Q(comparador_nonce_synth_1_11_) );
	DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_bF_buf39), .D(_933__12_), .Q(comparador_nonce_synth_1_12_) );
	DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_bF_buf38), .D(_933__13_), .Q(comparador_nonce_synth_1_13_) );
	DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_bF_buf37), .D(_933__14_), .Q(comparador_nonce_synth_1_14_) );
	DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_bF_buf36), .D(_933__15_), .Q(comparador_nonce_synth_1_15_) );
	DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_bF_buf35), .D(_933__16_), .Q(comparador_nonce_synth_1_16_) );
	DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_bF_buf34), .D(_933__17_), .Q(comparador_nonce_synth_1_17_) );
	DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_bF_buf33), .D(_933__18_), .Q(comparador_nonce_synth_1_18_) );
	DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_bF_buf32), .D(_933__19_), .Q(comparador_nonce_synth_1_19_) );
	DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_bF_buf31), .D(_933__20_), .Q(comparador_nonce_synth_1_20_) );
	DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_bF_buf30), .D(_933__21_), .Q(comparador_nonce_synth_1_21_) );
	DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_bF_buf29), .D(_933__22_), .Q(comparador_nonce_synth_1_22_) );
	DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_bF_buf28), .D(_933__23_), .Q(comparador_nonce_synth_1_23_) );
	DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_bF_buf27), .D(_933__24_), .Q(comparador_nonce_synth_1_24_) );
	DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_bF_buf26), .D(_933__25_), .Q(comparador_nonce_synth_1_25_) );
	DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_bF_buf25), .D(_933__26_), .Q(comparador_nonce_synth_1_26_) );
	DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_bF_buf24), .D(_933__27_), .Q(comparador_nonce_synth_1_27_) );
	DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_bF_buf23), .D(_933__28_), .Q(comparador_nonce_synth_1_28_) );
	DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_bF_buf22), .D(_933__29_), .Q(comparador_nonce_synth_1_29_) );
	DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_bF_buf21), .D(_933__30_), .Q(comparador_nonce_synth_1_30_) );
	DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_bF_buf20), .D(_933__31_), .Q(comparador_nonce_synth_1_31_) );
	DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_bF_buf19), .D(_928__0_), .Q(micro_hash_synth_a_0_) );
	DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_bF_buf18), .D(_928__1_), .Q(micro_hash_synth_a_1_) );
	DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_bF_buf17), .D(_928__2_), .Q(micro_hash_synth_a_2_) );
	DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_bF_buf16), .D(_928__3_), .Q(micro_hash_synth_a_3_) );
	DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_bF_buf15), .D(_928__4_), .Q(micro_hash_synth_a_4_) );
	DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_bF_buf14), .D(_928__5_), .Q(micro_hash_synth_a_5_) );
	DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_bF_buf13), .D(_928__6_), .Q(micro_hash_synth_a_6_) );
	DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_bF_buf12), .D(_928__7_), .Q(micro_hash_synth_a_7_) );
	DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_bF_buf11), .D(_929__0_), .Q(micro_hash_synth_b_0_) );
	DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_bF_buf10), .D(_929__1_), .Q(micro_hash_synth_b_1_) );
	DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_bF_buf9), .D(_929__2_), .Q(micro_hash_synth_b_2_) );
	DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_bF_buf8), .D(_929__3_), .Q(micro_hash_synth_b_3_) );
	DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_bF_buf7), .D(_929__4_), .Q(micro_hash_synth_b_4_) );
	DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_bF_buf6), .D(_929__5_), .Q(micro_hash_synth_b_5_) );
	DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_bF_buf5), .D(_929__6_), .Q(micro_hash_synth_b_6_) );
	DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_bF_buf4), .D(_929__7_), .Q(micro_hash_synth_b_7_) );
	DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_bF_buf3), .D(_930__0_), .Q(micro_hash_synth_c_0_) );
	DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_bF_buf2), .D(_930__1_), .Q(micro_hash_synth_c_1_) );
	DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_bF_buf1), .D(_930__2_), .Q(micro_hash_synth_c_2_) );
	DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_bF_buf0), .D(_930__3_), .Q(micro_hash_synth_c_3_) );
	DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_bF_buf76), .D(_930__4_), .Q(micro_hash_synth_c_4_) );
	DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_bF_buf75), .D(_930__5_), .Q(micro_hash_synth_c_5_) );
	DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_bF_buf74), .D(_930__6_), .Q(micro_hash_synth_c_6_) );
	DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_bF_buf73), .D(_930__7_), .Q(micro_hash_synth_c_7_) );
	DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_bF_buf72), .D(_932__0_), .Q(micro_hash_synth_k_0_) );
	DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_bF_buf71), .D(_932__1_), .Q(micro_hash_synth_k_1_) );
	DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_bF_buf70), .D(_932__2_), .Q(micro_hash_synth_k_2_) );
	DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_bF_buf69), .D(_932__3_), .Q(micro_hash_synth_k_3_) );
	DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_bF_buf68), .D(_932__4_), .Q(micro_hash_synth_k_4_) );
	DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_bF_buf67), .D(_932__5_), .Q(micro_hash_synth_k_5_) );
	DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_bF_buf66), .D(_932__6_), .Q(micro_hash_synth_k_6_) );
	DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_bF_buf65), .D(_932__7_), .Q(micro_hash_synth_k_7_) );
	DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_bF_buf64), .D(_934__0_), .Q(micro_hash_synth_x_0_) );
	DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_bF_buf63), .D(_934__1_), .Q(micro_hash_synth_x_1_) );
	DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_bF_buf62), .D(_934__2_), .Q(micro_hash_synth_x_2_) );
	DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_bF_buf61), .D(_934__3_), .Q(micro_hash_synth_x_3_) );
	DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_bF_buf60), .D(_934__4_), .Q(micro_hash_synth_x_4_) );
	DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_bF_buf59), .D(_934__5_), .Q(micro_hash_synth_x_5_) );
	DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_bF_buf58), .D(_934__6_), .Q(micro_hash_synth_x_6_) );
	DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_bF_buf57), .D(_934__7_), .Q(micro_hash_synth_x_7_) );
	DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_bF_buf56), .D(_1002_), .Q(micro_hash_synth_W_18__0_) );
	DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_bF_buf55), .D(_1004_), .Q(micro_hash_synth_W_18__1_) );
	DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_bF_buf54), .D(_1005_), .Q(micro_hash_synth_W_18__2_) );
	DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_bF_buf53), .D(_1006_), .Q(micro_hash_synth_W_18__3_) );
	DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_bF_buf52), .D(_1007_), .Q(micro_hash_synth_W_18__4_) );
	DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_bF_buf51), .D(_1008_), .Q(micro_hash_synth_W_18__5_) );
	DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_bF_buf50), .D(_1009_), .Q(micro_hash_synth_W_18__6_) );
	DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_bF_buf49), .D(_1010_), .Q(micro_hash_synth_W_18__7_) );
	DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_bF_buf48), .D(_1037_), .Q(micro_hash_synth_W_17__0_) );
	DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_bF_buf47), .D(_1038_), .Q(micro_hash_synth_W_17__1_) );
	DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_bF_buf46), .D(_1039_), .Q(micro_hash_synth_W_17__2_) );
	DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_bF_buf45), .D(_1040_), .Q(micro_hash_synth_W_17__3_) );
	DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_bF_buf44), .D(_1041_), .Q(micro_hash_synth_W_17__4_) );
	DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_bF_buf43), .D(_1042_), .Q(micro_hash_synth_W_17__5_) );
	DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_bF_buf42), .D(_1043_), .Q(micro_hash_synth_W_17__6_) );
	DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_bF_buf41), .D(_1044_), .Q(micro_hash_synth_W_17__7_) );
	DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_bF_buf40), .D(_1061_), .Q(micro_hash_synth_W_16__0_) );
	DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_bF_buf39), .D(_1062_), .Q(micro_hash_synth_W_16__1_) );
	DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_bF_buf38), .D(_1063_), .Q(micro_hash_synth_W_16__2_) );
	DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_bF_buf37), .D(_1064_), .Q(micro_hash_synth_W_16__3_) );
	DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_bF_buf36), .D(_1065_), .Q(micro_hash_synth_W_16__4_) );
	DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_bF_buf35), .D(_1066_), .Q(micro_hash_synth_W_16__5_) );
	DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_bF_buf34), .D(_1067_), .Q(micro_hash_synth_W_16__6_) );
	DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_bF_buf33), .D(_1068_), .Q(micro_hash_synth_W_16__7_) );
	DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_bF_buf32), .D(_977_), .Q(micro_hash_synth_W_15__0_) );
	DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_bF_buf31), .D(_978_), .Q(micro_hash_synth_W_15__1_) );
	DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_bF_buf30), .D(_979_), .Q(micro_hash_synth_W_15__2_) );
	DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_bF_buf29), .D(_980_), .Q(micro_hash_synth_W_15__3_) );
	DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_bF_buf28), .D(_981_), .Q(micro_hash_synth_W_15__4_) );
	DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_bF_buf27), .D(_982_), .Q(micro_hash_synth_W_15__5_) );
	DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_bF_buf26), .D(_983_), .Q(micro_hash_synth_W_15__6_) );
	DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_bF_buf25), .D(_984_), .Q(micro_hash_synth_W_15__7_) );
	DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_bF_buf24), .D(_1028_), .Q(micro_hash_synth_W_14__0_) );
	DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_bF_buf23), .D(_1029_), .Q(micro_hash_synth_W_14__1_) );
	DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_bF_buf22), .D(_1030_), .Q(micro_hash_synth_W_14__2_) );
	DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_bF_buf21), .D(_1031_), .Q(micro_hash_synth_W_14__3_) );
	DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_bF_buf20), .D(_1032_), .Q(micro_hash_synth_W_14__4_) );
	DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_bF_buf19), .D(_1033_), .Q(micro_hash_synth_W_14__5_) );
	DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_bF_buf18), .D(_1034_), .Q(micro_hash_synth_W_14__6_) );
	DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_bF_buf17), .D(_1036_), .Q(micro_hash_synth_W_14__7_) );
	DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_bF_buf16), .D(_1053_), .Q(micro_hash_synth_W_13__0_) );
	DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_bF_buf15), .D(_1054_), .Q(micro_hash_synth_W_13__1_) );
	DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_bF_buf14), .D(_1055_), .Q(micro_hash_synth_W_13__2_) );
	DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_bF_buf13), .D(_1056_), .Q(micro_hash_synth_W_13__3_) );
	DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_bF_buf12), .D(_1057_), .Q(micro_hash_synth_W_13__4_) );
	DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_bF_buf11), .D(_1058_), .Q(micro_hash_synth_W_13__5_) );
	DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_bF_buf10), .D(_1059_), .Q(micro_hash_synth_W_13__6_) );
	DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_bF_buf9), .D(_1060_), .Q(micro_hash_synth_W_13__7_) );
	DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_bF_buf8), .D(_1011_), .Q(micro_hash_synth_W_12__0_) );
	DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_bF_buf7), .D(_1012_), .Q(micro_hash_synth_W_12__1_) );
	DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_bF_buf6), .D(_1013_), .Q(micro_hash_synth_W_12__2_) );
	DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_bF_buf5), .D(_1014_), .Q(micro_hash_synth_W_12__3_) );
	DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_bF_buf4), .D(_1015_), .Q(micro_hash_synth_W_12__4_) );
	DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_bF_buf3), .D(_1016_), .Q(micro_hash_synth_W_12__5_) );
	DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_bF_buf2), .D(_1017_), .Q(micro_hash_synth_W_12__6_) );
	DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_bF_buf1), .D(_1018_), .Q(micro_hash_synth_W_12__7_) );
	DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_bF_buf0), .D(_1132_), .Q(micro_hash_synth_W_11__0_) );
	DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_bF_buf76), .D(_1133_), .Q(micro_hash_synth_W_11__1_) );
	DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_bF_buf75), .D(_1134_), .Q(micro_hash_synth_W_11__2_) );
	DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_bF_buf74), .D(_1135_), .Q(micro_hash_synth_W_11__3_) );
	DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_bF_buf73), .D(_1137_), .Q(micro_hash_synth_W_11__4_) );
	DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_bF_buf72), .D(_1138_), .Q(micro_hash_synth_W_11__5_) );
	DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_bF_buf71), .D(_1139_), .Q(micro_hash_synth_W_11__6_) );
	DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_bF_buf70), .D(_1140_), .Q(micro_hash_synth_W_11__7_) );
	DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_bF_buf69), .D(_1069_), .Q(micro_hash_synth_W_10__0_) );
	DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_bF_buf68), .D(_1070_), .Q(micro_hash_synth_W_10__1_) );
	DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_bF_buf67), .D(_1071_), .Q(micro_hash_synth_W_10__2_) );
	DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_bF_buf66), .D(_1072_), .Q(micro_hash_synth_W_10__3_) );
	DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_bF_buf65), .D(_1073_), .Q(micro_hash_synth_W_10__4_) );
	DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_bF_buf64), .D(_1074_), .Q(micro_hash_synth_W_10__5_) );
	DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_bF_buf63), .D(_1075_), .Q(micro_hash_synth_W_10__6_) );
	DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_bF_buf62), .D(_1076_), .Q(micro_hash_synth_W_10__7_) );
	DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_bF_buf61), .D(_1147_), .Q(micro_hash_synth_W_9__0_) );
	DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_bF_buf60), .D(_1158_), .Q(micro_hash_synth_W_9__1_) );
	DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_bF_buf59), .D(_1169_), .Q(micro_hash_synth_W_9__2_) );
	DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_bF_buf58), .D(_1176_), .Q(micro_hash_synth_W_9__3_) );
	DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_bF_buf57), .D(_1177_), .Q(micro_hash_synth_W_9__4_) );
	DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_bF_buf56), .D(_1178_), .Q(micro_hash_synth_W_9__5_) );
	DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_bF_buf55), .D(_1179_), .Q(micro_hash_synth_W_9__6_) );
	DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_bF_buf54), .D(_1180_), .Q(micro_hash_synth_W_9__7_) );
	DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_bF_buf53), .D(_1159_), .Q(micro_hash_synth_W_8__0_) );
	DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_bF_buf52), .D(_1160_), .Q(micro_hash_synth_W_8__1_) );
	DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_bF_buf51), .D(_1161_), .Q(micro_hash_synth_W_8__2_) );
	DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_bF_buf50), .D(_1162_), .Q(micro_hash_synth_W_8__3_) );
	DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_bF_buf49), .D(_1163_), .Q(micro_hash_synth_W_8__4_) );
	DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_bF_buf48), .D(_1164_), .Q(micro_hash_synth_W_8__5_) );
	DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_bF_buf47), .D(_1165_), .Q(micro_hash_synth_W_8__6_) );
	DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_bF_buf46), .D(_1166_), .Q(micro_hash_synth_W_8__7_) );
	DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_bF_buf45), .D(_1020_), .Q(micro_hash_synth_W_7__0_) );
	DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_bF_buf44), .D(_1021_), .Q(micro_hash_synth_W_7__1_) );
	DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_bF_buf43), .D(_1022_), .Q(micro_hash_synth_W_7__2_) );
	DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_bF_buf42), .D(_1023_), .Q(micro_hash_synth_W_7__3_) );
	DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_bF_buf41), .D(_1024_), .Q(micro_hash_synth_W_7__4_) );
	DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_bF_buf40), .D(_1025_), .Q(micro_hash_synth_W_7__5_) );
	DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_bF_buf39), .D(_1026_), .Q(micro_hash_synth_W_7__6_) );
	DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_bF_buf38), .D(_1027_), .Q(micro_hash_synth_W_7__7_) );
	DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_bF_buf37), .D(_968_), .Q(micro_hash_synth_W_6__0_) );
	DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_bF_buf36), .D(_969_), .Q(micro_hash_synth_W_6__1_) );
	DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_bF_buf35), .D(_970_), .Q(micro_hash_synth_W_6__2_) );
	DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_bF_buf34), .D(_972_), .Q(micro_hash_synth_W_6__3_) );
	DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_bF_buf33), .D(_973_), .Q(micro_hash_synth_W_6__4_) );
	DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_bF_buf32), .D(_974_), .Q(micro_hash_synth_W_6__5_) );
	DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_bF_buf31), .D(_975_), .Q(micro_hash_synth_W_6__6_) );
	DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_bF_buf30), .D(_976_), .Q(micro_hash_synth_W_6__7_) );
	DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_bF_buf29), .D(_1181_), .Q(micro_hash_synth_W_5__0_) );
	DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_bF_buf28), .D(_1182_), .Q(micro_hash_synth_W_5__1_) );
	DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_bF_buf27), .D(_1183_), .Q(micro_hash_synth_W_5__2_) );
	DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_bF_buf26), .D(_1184_), .Q(micro_hash_synth_W_5__3_) );
	DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_bF_buf25), .D(_1185_), .Q(micro_hash_synth_W_5__4_) );
	DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_bF_buf24), .D(_1186_), .Q(micro_hash_synth_W_5__5_) );
	DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_bF_buf23), .D(_1187_), .Q(micro_hash_synth_W_5__6_) );
	DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_bF_buf22), .D(_1189_), .Q(micro_hash_synth_W_5__7_) );
	DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_bF_buf21), .D(_1123_), .Q(micro_hash_synth_W_4__0_) );
	DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_bF_buf20), .D(_1124_), .Q(micro_hash_synth_W_4__1_) );
	DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_bF_buf19), .D(_1126_), .Q(micro_hash_synth_W_4__2_) );
	DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_bF_buf18), .D(_1127_), .Q(micro_hash_synth_W_4__3_) );
	DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_bF_buf17), .D(_1128_), .Q(micro_hash_synth_W_4__4_) );
	DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_bF_buf16), .D(_1129_), .Q(micro_hash_synth_W_4__5_) );
	DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_bF_buf15), .D(_1130_), .Q(micro_hash_synth_W_4__6_) );
	DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_bF_buf14), .D(_1131_), .Q(micro_hash_synth_W_4__7_) );
	DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_bF_buf13), .D(_1150_), .Q(micro_hash_synth_W_23__0_) );
	DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_bF_buf12), .D(_1151_), .Q(micro_hash_synth_W_23__1_) );
	DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_bF_buf11), .D(_1152_), .Q(micro_hash_synth_W_23__2_) );
	DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_bF_buf10), .D(_1153_), .Q(micro_hash_synth_W_23__3_) );
	DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_bF_buf9), .D(_1154_), .Q(micro_hash_synth_W_23__4_) );
	DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_bF_buf8), .D(_1155_), .Q(micro_hash_synth_W_23__5_) );
	DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_bF_buf7), .D(_1156_), .Q(micro_hash_synth_W_23__6_) );
	DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_bF_buf6), .D(_1157_), .Q(micro_hash_synth_W_23__7_) );
	DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_bF_buf5), .D(_1141_), .Q(micro_hash_synth_W_24__0_) );
	DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_bF_buf4), .D(_1142_), .Q(micro_hash_synth_W_24__1_) );
	DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_bF_buf3), .D(_1143_), .Q(micro_hash_synth_W_24__2_) );
	DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_bF_buf2), .D(_1144_), .Q(micro_hash_synth_W_24__3_) );
	DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_bF_buf1), .D(_1145_), .Q(micro_hash_synth_W_24__4_) );
	DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_bF_buf0), .D(_1146_), .Q(micro_hash_synth_W_24__5_) );
	DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_bF_buf76), .D(_1148_), .Q(micro_hash_synth_W_24__6_) );
	DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_bF_buf75), .D(_1149_), .Q(micro_hash_synth_W_24__7_) );
	DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_bF_buf74), .D(_941_), .Q(micro_hash_synth_W_25__0_) );
	DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_bF_buf73), .D(_950_), .Q(micro_hash_synth_W_25__1_) );
	DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_bF_buf72), .D(_955_), .Q(micro_hash_synth_W_25__2_) );
	DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_bF_buf71), .D(_971_), .Q(micro_hash_synth_W_25__3_) );
	DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_bF_buf70), .D(_987_), .Q(micro_hash_synth_W_25__4_) );
	DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_bF_buf69), .D(_1003_), .Q(micro_hash_synth_W_25__5_) );
	DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_bF_buf68), .D(_1019_), .Q(micro_hash_synth_W_25__6_) );
	DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_bF_buf67), .D(_1035_), .Q(micro_hash_synth_W_25__7_) );
	DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_bF_buf66), .D(_1188_), .Q(micro_hash_synth_W_26__0_) );
	DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_bF_buf65), .D(_1190_), .Q(micro_hash_synth_W_26__1_) );
	DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_bF_buf64), .D(_935_), .Q(micro_hash_synth_W_26__2_) );
	DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_bF_buf63), .D(_936_), .Q(micro_hash_synth_W_26__3_) );
	DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_bF_buf62), .D(_937_), .Q(micro_hash_synth_W_26__4_) );
	DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_bF_buf61), .D(_938_), .Q(micro_hash_synth_W_26__5_) );
	DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_bF_buf60), .D(_939_), .Q(micro_hash_synth_W_26__6_) );
	DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_bF_buf59), .D(_940_), .Q(micro_hash_synth_W_26__7_) );
	DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_bF_buf58), .D(_1115_), .Q(micro_hash_synth_W_3__0_) );
	DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_bF_buf57), .D(_1116_), .Q(micro_hash_synth_W_3__1_) );
	DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_bF_buf56), .D(_1117_), .Q(micro_hash_synth_W_3__2_) );
	DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_bF_buf55), .D(_1118_), .Q(micro_hash_synth_W_3__3_) );
	DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_bF_buf54), .D(_1119_), .Q(micro_hash_synth_W_3__4_) );
	DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_bF_buf53), .D(_1120_), .Q(micro_hash_synth_W_3__5_) );
	DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_bF_buf52), .D(_1121_), .Q(micro_hash_synth_W_3__6_) );
	DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_bF_buf51), .D(_1122_), .Q(micro_hash_synth_W_3__7_) );
	DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_bF_buf50), .D(_1109_), .Q(micro_hash_synth_W_27__0_) );
	DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_bF_buf49), .D(_1110_), .Q(micro_hash_synth_W_27__1_) );
	DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_bF_buf48), .D(_1111_), .Q(micro_hash_synth_W_27__2_) );
	DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_bF_buf47), .D(_1112_), .Q(micro_hash_synth_W_27__3_) );
	DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_bF_buf46), .D(_1113_), .Q(micro_hash_synth_W_27__4_) );
	DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_bF_buf45), .D(_1114_), .Q(micro_hash_synth_W_27__5_) );
	DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_bF_buf44), .D(_1125_), .Q(micro_hash_synth_W_27__6_) );
	DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_bF_buf43), .D(_1136_), .Q(micro_hash_synth_W_27__7_) );
	DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_bF_buf42), .D(_1077_), .Q(micro_hash_synth_W_28__0_) );
	DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_bF_buf41), .D(_1078_), .Q(micro_hash_synth_W_28__1_) );
	DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_bF_buf40), .D(_1079_), .Q(micro_hash_synth_W_28__2_) );
	DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_bF_buf39), .D(_1080_), .Q(micro_hash_synth_W_28__3_) );
	DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_bF_buf38), .D(_1081_), .Q(micro_hash_synth_W_28__4_) );
	DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_bF_buf37), .D(_1082_), .Q(micro_hash_synth_W_28__5_) );
	DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_bF_buf36), .D(_1083_), .Q(micro_hash_synth_W_28__6_) );
	DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_bF_buf35), .D(_1084_), .Q(micro_hash_synth_W_28__7_) );
	DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_bF_buf34), .D(_1085_), .Q(micro_hash_synth_W_29__0_) );
	DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_bF_buf33), .D(_1086_), .Q(micro_hash_synth_W_29__1_) );
	DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_bF_buf32), .D(_1087_), .Q(micro_hash_synth_W_29__2_) );
	DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_bF_buf31), .D(_1088_), .Q(micro_hash_synth_W_29__3_) );
	DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_bF_buf30), .D(_1089_), .Q(micro_hash_synth_W_29__4_) );
	DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_bF_buf29), .D(_1090_), .Q(micro_hash_synth_W_29__5_) );
	DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_bF_buf28), .D(_1091_), .Q(micro_hash_synth_W_29__6_) );
	DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_bF_buf27), .D(_1092_), .Q(micro_hash_synth_W_29__7_) );
	DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_bF_buf26), .D(_1093_), .Q(micro_hash_synth_W_30__0_) );
	DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_bF_buf25), .D(_1094_), .Q(micro_hash_synth_W_30__1_) );
	DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_bF_buf24), .D(_1095_), .Q(micro_hash_synth_W_30__2_) );
	DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_bF_buf23), .D(_1096_), .Q(micro_hash_synth_W_30__3_) );
	DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_bF_buf22), .D(_1097_), .Q(micro_hash_synth_W_30__4_) );
	DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_bF_buf21), .D(_1098_), .Q(micro_hash_synth_W_30__5_) );
	DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_bF_buf20), .D(_1099_), .Q(micro_hash_synth_W_30__6_) );
	DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_bF_buf19), .D(_1100_), .Q(micro_hash_synth_W_30__7_) );
	DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_bF_buf18), .D(_1101_), .Q(micro_hash_synth_W_31__0_) );
	DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_bF_buf17), .D(_1102_), .Q(micro_hash_synth_W_31__1_) );
	DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_bF_buf16), .D(_1103_), .Q(micro_hash_synth_W_31__2_) );
	DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_bF_buf15), .D(_1104_), .Q(micro_hash_synth_W_31__3_) );
	DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_bF_buf14), .D(_1105_), .Q(micro_hash_synth_W_31__4_) );
	DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_bF_buf13), .D(_1106_), .Q(micro_hash_synth_W_31__5_) );
	DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_bF_buf12), .D(_1107_), .Q(micro_hash_synth_W_31__6_) );
	DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_bF_buf11), .D(_1108_), .Q(micro_hash_synth_W_31__7_) );
	DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_bF_buf10), .D(_994_), .Q(micro_hash_synth_W_1__0_) );
	DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_bF_buf9), .D(_995_), .Q(micro_hash_synth_W_1__1_) );
	DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_bF_buf8), .D(_996_), .Q(micro_hash_synth_W_1__2_) );
	DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_bF_buf7), .D(_997_), .Q(micro_hash_synth_W_1__3_) );
	DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_bF_buf6), .D(_998_), .Q(micro_hash_synth_W_1__4_) );
	DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_bF_buf5), .D(_999_), .Q(micro_hash_synth_W_1__5_) );
	DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_bF_buf4), .D(_1000_), .Q(micro_hash_synth_W_1__6_) );
	DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_bF_buf3), .D(_1001_), .Q(micro_hash_synth_W_1__7_) );
	DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_bF_buf2), .D(_1045_), .Q(micro_hash_synth_W_2__0_) );
	DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_bF_buf1), .D(_1046_), .Q(micro_hash_synth_W_2__1_) );
	DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_bF_buf0), .D(_1047_), .Q(micro_hash_synth_W_2__2_) );
	DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_bF_buf76), .D(_1048_), .Q(micro_hash_synth_W_2__3_) );
	DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_bF_buf75), .D(_1049_), .Q(micro_hash_synth_W_2__4_) );
	DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_bF_buf74), .D(_1050_), .Q(micro_hash_synth_W_2__5_) );
	DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_bF_buf73), .D(_1051_), .Q(micro_hash_synth_W_2__6_) );
	DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_bF_buf72), .D(_1052_), .Q(micro_hash_synth_W_2__7_) );
	INVX8 INVX8_5 ( .A(reset_L_bF_buf10), .Y(_2618_) );
	INVX1 INVX1_655 ( .A(num_entradas[1]), .Y(_2619_) );
	INVX1 INVX1_656 ( .A(num_entradas[0]), .Y(_2620_) );
	OAI22X1 OAI22X1_269 ( .A(_2619_), .B(RAM_rd_ptr_1_), .C(_2620_), .D(RAM_rd_ptr_0_), .Y(_2621_) );
	INVX1 INVX1_657 ( .A(comparador_valid_bF_buf2), .Y(_2622_) );
	AOI21X1 AOI21X1_446 ( .A(RAM_rd_ptr_1_), .B(_2619_), .C(_2622_), .Y(_2623_) );
	AOI21X1 AOI21X1_447 ( .A(RAM_rd_ptr_0_), .B(_2620_), .C(_1__bF_buf4), .Y(_2624_) );
	OAI21X1 OAI21X1_661 ( .A(_2621_), .B(_2624_), .C(_2623_), .Y(_2625_) );
	NAND2X1 NAND2X1_264 ( .A(_3__0_), .B(_2625__bF_buf6), .Y(_2626_) );
	INVX1 INVX1_658 ( .A(RAM_rd_ptr_1_), .Y(_2627_) );
	INVX1 INVX1_659 ( .A(RAM_rd_ptr_0_), .Y(_2628_) );
	AOI22X1 AOI22X1_64 ( .A(_2627_), .B(num_entradas[1]), .C(num_entradas[0]), .D(_2628_), .Y(_2629_) );
	OAI21X1 OAI21X1_662 ( .A(_2627_), .B(num_entradas[1]), .C(comparador_valid_bF_buf1), .Y(_2630_) );
	INVX1 INVX1_660 ( .A(_1__bF_buf3), .Y(_2631_) );
	OAI21X1 OAI21X1_663 ( .A(_2628_), .B(num_entradas[0]), .C(_2631_), .Y(_2632_) );
	AOI21X1 AOI21X1_448 ( .A(_2632_), .B(_2629_), .C(_2630_), .Y(_2633_) );
	NAND2X1 NAND2X1_265 ( .A(comparador_nonce_synth_valido_0_), .B(_2633__bF_buf6), .Y(_2634_) );
	AOI21X1 AOI21X1_449 ( .A(_2626_), .B(_2634_), .C(_2618__bF_buf6), .Y(_2616__0_) );
	NAND2X1 NAND2X1_266 ( .A(_3__1_), .B(_2625__bF_buf5), .Y(_2635_) );
	NAND2X1 NAND2X1_267 ( .A(comparador_nonce_synth_valido_1_), .B(_2633__bF_buf5), .Y(_2636_) );
	AOI21X1 AOI21X1_450 ( .A(_2635_), .B(_2636_), .C(_2618__bF_buf5), .Y(_2616__1_) );
	NAND2X1 NAND2X1_268 ( .A(_3__2_), .B(_2625__bF_buf4), .Y(_2637_) );
	NAND2X1 NAND2X1_269 ( .A(comparador_nonce_synth_valido_2_), .B(_2633__bF_buf4), .Y(_2638_) );
	AOI21X1 AOI21X1_451 ( .A(_2637_), .B(_2638_), .C(_2618__bF_buf4), .Y(_2616__2_) );
	NAND2X1 NAND2X1_270 ( .A(_3__3_), .B(_2625__bF_buf3), .Y(_2639_) );
	NAND2X1 NAND2X1_271 ( .A(comparador_nonce_synth_valido_3_), .B(_2633__bF_buf3), .Y(_2640_) );
	AOI21X1 AOI21X1_452 ( .A(_2639_), .B(_2640_), .C(_2618__bF_buf3), .Y(_2616__3_) );
	NAND2X1 NAND2X1_272 ( .A(_3__4_), .B(_2625__bF_buf2), .Y(_2641_) );
	NAND2X1 NAND2X1_273 ( .A(comparador_nonce_synth_valido_4_), .B(_2633__bF_buf2), .Y(_2642_) );
	AOI21X1 AOI21X1_453 ( .A(_2641_), .B(_2642_), .C(_2618__bF_buf2), .Y(_2616__4_) );
	NAND2X1 NAND2X1_274 ( .A(_3__5_), .B(_2625__bF_buf1), .Y(_2643_) );
	NAND2X1 NAND2X1_275 ( .A(comparador_nonce_synth_valido_5_), .B(_2633__bF_buf1), .Y(_2644_) );
	AOI21X1 AOI21X1_454 ( .A(_2643_), .B(_2644_), .C(_2618__bF_buf1), .Y(_2616__5_) );
	NAND2X1 NAND2X1_276 ( .A(_3__6_), .B(_2625__bF_buf0), .Y(_2645_) );
	NAND2X1 NAND2X1_277 ( .A(comparador_nonce_synth_valido_6_), .B(_2633__bF_buf0), .Y(_2646_) );
	AOI21X1 AOI21X1_455 ( .A(_2645_), .B(_2646_), .C(_2618__bF_buf0), .Y(_2616__6_) );
	NAND2X1 NAND2X1_278 ( .A(_3__7_), .B(_2625__bF_buf6), .Y(_2647_) );
	NAND2X1 NAND2X1_279 ( .A(comparador_nonce_synth_valido_7_), .B(_2633__bF_buf6), .Y(_2648_) );
	AOI21X1 AOI21X1_456 ( .A(_2647_), .B(_2648_), .C(_2618__bF_buf6), .Y(_2616__7_) );
	NAND2X1 NAND2X1_280 ( .A(_3__8_), .B(_2625__bF_buf5), .Y(_2649_) );
	NAND2X1 NAND2X1_281 ( .A(comparador_nonce_synth_valido_8_), .B(_2633__bF_buf5), .Y(_2650_) );
	AOI21X1 AOI21X1_457 ( .A(_2649_), .B(_2650_), .C(_2618__bF_buf5), .Y(_2616__8_) );
	NAND2X1 NAND2X1_282 ( .A(_3__9_), .B(_2625__bF_buf4), .Y(_2651_) );
	NAND2X1 NAND2X1_283 ( .A(comparador_nonce_synth_valido_9_), .B(_2633__bF_buf4), .Y(_2652_) );
	AOI21X1 AOI21X1_458 ( .A(_2651_), .B(_2652_), .C(_2618__bF_buf4), .Y(_2616__9_) );
	NAND2X1 NAND2X1_284 ( .A(_3__10_), .B(_2625__bF_buf3), .Y(_2653_) );
	NAND2X1 NAND2X1_285 ( .A(comparador_nonce_synth_valido_10_), .B(_2633__bF_buf3), .Y(_2654_) );
	AOI21X1 AOI21X1_459 ( .A(_2653_), .B(_2654_), .C(_2618__bF_buf3), .Y(_2616__10_) );
	NAND2X1 NAND2X1_286 ( .A(_3__11_), .B(_2625__bF_buf2), .Y(_2655_) );
	NAND2X1 NAND2X1_287 ( .A(comparador_nonce_synth_valido_11_), .B(_2633__bF_buf2), .Y(_2656_) );
	AOI21X1 AOI21X1_460 ( .A(_2655_), .B(_2656_), .C(_2618__bF_buf2), .Y(_2616__11_) );
	NAND2X1 NAND2X1_288 ( .A(_3__12_), .B(_2625__bF_buf1), .Y(_2657_) );
	NAND2X1 NAND2X1_289 ( .A(comparador_nonce_synth_valido_12_), .B(_2633__bF_buf1), .Y(_2658_) );
	AOI21X1 AOI21X1_461 ( .A(_2657_), .B(_2658_), .C(_2618__bF_buf1), .Y(_2616__12_) );
	NAND2X1 NAND2X1_290 ( .A(_3__13_), .B(_2625__bF_buf0), .Y(_2659_) );
	NAND2X1 NAND2X1_291 ( .A(comparador_nonce_synth_valido_13_), .B(_2633__bF_buf0), .Y(_2660_) );
	AOI21X1 AOI21X1_462 ( .A(_2659_), .B(_2660_), .C(_2618__bF_buf0), .Y(_2616__13_) );
	NAND2X1 NAND2X1_292 ( .A(_3__14_), .B(_2625__bF_buf6), .Y(_2661_) );
	NAND2X1 NAND2X1_293 ( .A(comparador_nonce_synth_valido_14_), .B(_2633__bF_buf6), .Y(_2662_) );
	AOI21X1 AOI21X1_463 ( .A(_2661_), .B(_2662_), .C(_2618__bF_buf6), .Y(_2616__14_) );
	NAND2X1 NAND2X1_294 ( .A(_3__15_), .B(_2625__bF_buf5), .Y(_2663_) );
	NAND2X1 NAND2X1_295 ( .A(comparador_nonce_synth_valido_15_), .B(_2633__bF_buf5), .Y(_2664_) );
	AOI21X1 AOI21X1_464 ( .A(_2663_), .B(_2664_), .C(_2618__bF_buf5), .Y(_2616__15_) );
	NAND2X1 NAND2X1_296 ( .A(_3__16_), .B(_2625__bF_buf4), .Y(_2665_) );
	NAND2X1 NAND2X1_297 ( .A(comparador_nonce_synth_valido_16_), .B(_2633__bF_buf4), .Y(_2666_) );
	AOI21X1 AOI21X1_465 ( .A(_2665_), .B(_2666_), .C(_2618__bF_buf4), .Y(_2616__16_) );
	NAND2X1 NAND2X1_298 ( .A(_3__17_), .B(_2625__bF_buf3), .Y(_2667_) );
	NAND2X1 NAND2X1_299 ( .A(comparador_nonce_synth_valido_17_), .B(_2633__bF_buf3), .Y(_2668_) );
	AOI21X1 AOI21X1_466 ( .A(_2667_), .B(_2668_), .C(_2618__bF_buf3), .Y(_2616__17_) );
	NAND2X1 NAND2X1_300 ( .A(_3__18_), .B(_2625__bF_buf2), .Y(_2669_) );
	NAND2X1 NAND2X1_301 ( .A(comparador_nonce_synth_valido_18_), .B(_2633__bF_buf2), .Y(_2670_) );
	AOI21X1 AOI21X1_467 ( .A(_2669_), .B(_2670_), .C(_2618__bF_buf2), .Y(_2616__18_) );
	NAND2X1 NAND2X1_302 ( .A(_3__19_), .B(_2625__bF_buf1), .Y(_2671_) );
	NAND2X1 NAND2X1_303 ( .A(comparador_nonce_synth_valido_19_), .B(_2633__bF_buf1), .Y(_2672_) );
	AOI21X1 AOI21X1_468 ( .A(_2671_), .B(_2672_), .C(_2618__bF_buf1), .Y(_2616__19_) );
	NAND2X1 NAND2X1_304 ( .A(_3__20_), .B(_2625__bF_buf0), .Y(_2673_) );
	NAND2X1 NAND2X1_305 ( .A(comparador_nonce_synth_valido_20_), .B(_2633__bF_buf0), .Y(_2674_) );
	AOI21X1 AOI21X1_469 ( .A(_2673_), .B(_2674_), .C(_2618__bF_buf0), .Y(_2616__20_) );
	NAND2X1 NAND2X1_306 ( .A(_3__21_), .B(_2625__bF_buf6), .Y(_2675_) );
	NAND2X1 NAND2X1_307 ( .A(comparador_nonce_synth_valido_21_), .B(_2633__bF_buf6), .Y(_2676_) );
	AOI21X1 AOI21X1_470 ( .A(_2675_), .B(_2676_), .C(_2618__bF_buf6), .Y(_2616__21_) );
	NAND2X1 NAND2X1_308 ( .A(_3__22_), .B(_2625__bF_buf5), .Y(_2677_) );
	NAND2X1 NAND2X1_309 ( .A(comparador_nonce_synth_valido_22_), .B(_2633__bF_buf5), .Y(_2678_) );
	AOI21X1 AOI21X1_471 ( .A(_2677_), .B(_2678_), .C(_2618__bF_buf5), .Y(_2616__22_) );
	NAND2X1 NAND2X1_310 ( .A(_3__23_), .B(_2625__bF_buf4), .Y(_2679_) );
	NAND2X1 NAND2X1_311 ( .A(comparador_nonce_synth_valido_23_), .B(_2633__bF_buf4), .Y(_2680_) );
	AOI21X1 AOI21X1_472 ( .A(_2679_), .B(_2680_), .C(_2618__bF_buf4), .Y(_2616__23_) );
	NAND2X1 NAND2X1_312 ( .A(_3__24_), .B(_2625__bF_buf3), .Y(_2681_) );
	NAND2X1 NAND2X1_313 ( .A(comparador_nonce_synth_valido_24_), .B(_2633__bF_buf3), .Y(_2682_) );
	AOI21X1 AOI21X1_473 ( .A(_2681_), .B(_2682_), .C(_2618__bF_buf3), .Y(_2616__24_) );
	NAND2X1 NAND2X1_314 ( .A(_3__25_), .B(_2625__bF_buf2), .Y(_2683_) );
	NAND2X1 NAND2X1_315 ( .A(comparador_nonce_synth_valido_25_), .B(_2633__bF_buf2), .Y(_2684_) );
	AOI21X1 AOI21X1_474 ( .A(_2683_), .B(_2684_), .C(_2618__bF_buf2), .Y(_2616__25_) );
	NAND2X1 NAND2X1_316 ( .A(_3__26_), .B(_2625__bF_buf1), .Y(_2685_) );
	NAND2X1 NAND2X1_317 ( .A(comparador_nonce_synth_valido_26_), .B(_2633__bF_buf1), .Y(_2686_) );
	AOI21X1 AOI21X1_475 ( .A(_2685_), .B(_2686_), .C(_2618__bF_buf1), .Y(_2616__26_) );
	NAND2X1 NAND2X1_318 ( .A(_3__27_), .B(_2625__bF_buf0), .Y(_2687_) );
	NAND2X1 NAND2X1_319 ( .A(comparador_nonce_synth_valido_27_), .B(_2633__bF_buf0), .Y(_2688_) );
	AOI21X1 AOI21X1_476 ( .A(_2687_), .B(_2688_), .C(_2618__bF_buf0), .Y(_2616__27_) );
	NAND2X1 NAND2X1_320 ( .A(_3__28_), .B(_2625__bF_buf6), .Y(_2689_) );
	NAND2X1 NAND2X1_321 ( .A(comparador_nonce_synth_valido_28_), .B(_2633__bF_buf6), .Y(_2690_) );
	AOI21X1 AOI21X1_477 ( .A(_2689_), .B(_2690_), .C(_2618__bF_buf6), .Y(_2616__28_) );
	NAND2X1 NAND2X1_322 ( .A(_3__29_), .B(_2625__bF_buf5), .Y(_2691_) );
	NAND2X1 NAND2X1_323 ( .A(comparador_nonce_synth_valido_29_), .B(_2633__bF_buf5), .Y(_2692_) );
	AOI21X1 AOI21X1_478 ( .A(_2691_), .B(_2692_), .C(_2618__bF_buf5), .Y(_2616__29_) );
	NAND2X1 NAND2X1_324 ( .A(_3__30_), .B(_2625__bF_buf4), .Y(_2693_) );
	NAND2X1 NAND2X1_325 ( .A(comparador_nonce_synth_valido_30_), .B(_2633__bF_buf4), .Y(_2694_) );
	AOI21X1 AOI21X1_479 ( .A(_2693_), .B(_2694_), .C(_2618__bF_buf4), .Y(_2616__30_) );
	NAND2X1 NAND2X1_326 ( .A(_3__31_), .B(_2625__bF_buf3), .Y(_2695_) );
	NAND2X1 NAND2X1_327 ( .A(comparador_nonce_synth_valido_31_), .B(_2633__bF_buf3), .Y(_2696_) );
	AOI21X1 AOI21X1_480 ( .A(_2695_), .B(_2696_), .C(_2618__bF_buf3), .Y(_2616__31_) );
	NAND2X1 NAND2X1_328 ( .A(_0__0_), .B(_2625__bF_buf2), .Y(_2697_) );
	NAND2X1 NAND2X1_329 ( .A(bounty_synth_0_), .B(_2633__bF_buf2), .Y(_2698_) );
	AOI21X1 AOI21X1_481 ( .A(_2697_), .B(_2698_), .C(_2618__bF_buf2), .Y(_2614__0_) );
	NAND2X1 NAND2X1_330 ( .A(_0__1_), .B(_2625__bF_buf1), .Y(_2699_) );
	NAND2X1 NAND2X1_331 ( .A(bounty_synth_1_), .B(_2633__bF_buf1), .Y(_2700_) );
	AOI21X1 AOI21X1_482 ( .A(_2699_), .B(_2700_), .C(_2618__bF_buf1), .Y(_2614__1_) );
	NAND2X1 NAND2X1_332 ( .A(_0__2_), .B(_2625__bF_buf0), .Y(_2701_) );
	NAND2X1 NAND2X1_333 ( .A(bounty_synth_2_), .B(_2633__bF_buf0), .Y(_2702_) );
	AOI21X1 AOI21X1_483 ( .A(_2701_), .B(_2702_), .C(_2618__bF_buf0), .Y(_2614__2_) );
	NAND2X1 NAND2X1_334 ( .A(_0__3_), .B(_2625__bF_buf6), .Y(_2703_) );
	NAND2X1 NAND2X1_335 ( .A(bounty_synth_3_), .B(_2633__bF_buf6), .Y(_2704_) );
	AOI21X1 AOI21X1_484 ( .A(_2703_), .B(_2704_), .C(_2618__bF_buf6), .Y(_2614__3_) );
	NAND2X1 NAND2X1_336 ( .A(_0__4_), .B(_2625__bF_buf5), .Y(_2705_) );
	NAND2X1 NAND2X1_337 ( .A(bounty_synth_4_), .B(_2633__bF_buf5), .Y(_2706_) );
	AOI21X1 AOI21X1_485 ( .A(_2705_), .B(_2706_), .C(_2618__bF_buf5), .Y(_2614__4_) );
	NAND2X1 NAND2X1_338 ( .A(_0__5_), .B(_2625__bF_buf4), .Y(_2707_) );
	NAND2X1 NAND2X1_339 ( .A(bounty_synth_5_), .B(_2633__bF_buf4), .Y(_2708_) );
	AOI21X1 AOI21X1_486 ( .A(_2707_), .B(_2708_), .C(_2618__bF_buf4), .Y(_2614__5_) );
	NAND2X1 NAND2X1_340 ( .A(_0__6_), .B(_2625__bF_buf3), .Y(_2709_) );
	NAND2X1 NAND2X1_341 ( .A(bounty_synth_6_), .B(_2633__bF_buf3), .Y(_2710_) );
	AOI21X1 AOI21X1_487 ( .A(_2709_), .B(_2710_), .C(_2618__bF_buf3), .Y(_2614__6_) );
	NAND2X1 NAND2X1_342 ( .A(_0__7_), .B(_2625__bF_buf2), .Y(_2711_) );
	NAND2X1 NAND2X1_343 ( .A(bounty_synth_7_), .B(_2633__bF_buf2), .Y(_2712_) );
	AOI21X1 AOI21X1_488 ( .A(_2711_), .B(_2712_), .C(_2618__bF_buf2), .Y(_2614__7_) );
	NAND2X1 NAND2X1_344 ( .A(_0__8_), .B(_2625__bF_buf1), .Y(_2713_) );
	NAND2X1 NAND2X1_345 ( .A(bounty_synth_8_), .B(_2633__bF_buf1), .Y(_2714_) );
	AOI21X1 AOI21X1_489 ( .A(_2713_), .B(_2714_), .C(_2618__bF_buf1), .Y(_2614__8_) );
	NAND2X1 NAND2X1_346 ( .A(_0__9_), .B(_2625__bF_buf0), .Y(_2715_) );
	NAND2X1 NAND2X1_347 ( .A(bounty_synth_9_), .B(_2633__bF_buf0), .Y(_2716_) );
	AOI21X1 AOI21X1_490 ( .A(_2715_), .B(_2716_), .C(_2618__bF_buf0), .Y(_2614__9_) );
	NAND2X1 NAND2X1_348 ( .A(_0__10_), .B(_2625__bF_buf6), .Y(_2717_) );
	NAND2X1 NAND2X1_349 ( .A(bounty_synth_10_), .B(_2633__bF_buf6), .Y(_2718_) );
	AOI21X1 AOI21X1_491 ( .A(_2717_), .B(_2718_), .C(_2618__bF_buf6), .Y(_2614__10_) );
	NAND2X1 NAND2X1_350 ( .A(_0__11_), .B(_2625__bF_buf5), .Y(_2719_) );
	NAND2X1 NAND2X1_351 ( .A(bounty_synth_11_), .B(_2633__bF_buf5), .Y(_2720_) );
	AOI21X1 AOI21X1_492 ( .A(_2719_), .B(_2720_), .C(_2618__bF_buf5), .Y(_2614__11_) );
	NAND2X1 NAND2X1_352 ( .A(_0__12_), .B(_2625__bF_buf4), .Y(_2721_) );
	NAND2X1 NAND2X1_353 ( .A(bounty_synth_12_), .B(_2633__bF_buf4), .Y(_2722_) );
	AOI21X1 AOI21X1_493 ( .A(_2721_), .B(_2722_), .C(_2618__bF_buf4), .Y(_2614__12_) );
	NAND2X1 NAND2X1_354 ( .A(_0__13_), .B(_2625__bF_buf3), .Y(_2723_) );
	NAND2X1 NAND2X1_355 ( .A(bounty_synth_13_), .B(_2633__bF_buf3), .Y(_2724_) );
	AOI21X1 AOI21X1_494 ( .A(_2723_), .B(_2724_), .C(_2618__bF_buf3), .Y(_2614__13_) );
	NAND2X1 NAND2X1_356 ( .A(_0__14_), .B(_2625__bF_buf2), .Y(_2725_) );
	NAND2X1 NAND2X1_357 ( .A(bounty_synth_14_), .B(_2633__bF_buf2), .Y(_2726_) );
	AOI21X1 AOI21X1_495 ( .A(_2725_), .B(_2726_), .C(_2618__bF_buf2), .Y(_2614__14_) );
	NAND2X1 NAND2X1_358 ( .A(_0__15_), .B(_2625__bF_buf1), .Y(_2727_) );
	NAND2X1 NAND2X1_359 ( .A(bounty_synth_15_), .B(_2633__bF_buf1), .Y(_2728_) );
	AOI21X1 AOI21X1_496 ( .A(_2727_), .B(_2728_), .C(_2618__bF_buf1), .Y(_2614__15_) );
	NAND2X1 NAND2X1_360 ( .A(_0__16_), .B(_2625__bF_buf0), .Y(_2729_) );
	NAND2X1 NAND2X1_361 ( .A(bounty_synth_16_), .B(_2633__bF_buf0), .Y(_2730_) );
	AOI21X1 AOI21X1_497 ( .A(_2729_), .B(_2730_), .C(_2618__bF_buf0), .Y(_2614__16_) );
	NAND2X1 NAND2X1_362 ( .A(_0__17_), .B(_2625__bF_buf6), .Y(_2731_) );
	NAND2X1 NAND2X1_363 ( .A(bounty_synth_17_), .B(_2633__bF_buf6), .Y(_2732_) );
	AOI21X1 AOI21X1_498 ( .A(_2731_), .B(_2732_), .C(_2618__bF_buf6), .Y(_2614__17_) );
	NAND2X1 NAND2X1_364 ( .A(_0__18_), .B(_2625__bF_buf5), .Y(_2733_) );
	NAND2X1 NAND2X1_365 ( .A(bounty_synth_18_), .B(_2633__bF_buf5), .Y(_2734_) );
	AOI21X1 AOI21X1_499 ( .A(_2733_), .B(_2734_), .C(_2618__bF_buf5), .Y(_2614__18_) );
	NAND2X1 NAND2X1_366 ( .A(_0__19_), .B(_2625__bF_buf4), .Y(_2735_) );
	NAND2X1 NAND2X1_367 ( .A(bounty_synth_19_), .B(_2633__bF_buf4), .Y(_2736_) );
	AOI21X1 AOI21X1_500 ( .A(_2735_), .B(_2736_), .C(_2618__bF_buf4), .Y(_2614__19_) );
	NAND2X1 NAND2X1_368 ( .A(_0__20_), .B(_2625__bF_buf3), .Y(_2737_) );
	NAND2X1 NAND2X1_369 ( .A(bounty_synth_20_), .B(_2633__bF_buf3), .Y(_2738_) );
	AOI21X1 AOI21X1_501 ( .A(_2737_), .B(_2738_), .C(_2618__bF_buf3), .Y(_2614__20_) );
	NAND2X1 NAND2X1_370 ( .A(_0__21_), .B(_2625__bF_buf2), .Y(_2739_) );
	NAND2X1 NAND2X1_371 ( .A(bounty_synth_21_), .B(_2633__bF_buf2), .Y(_2740_) );
	AOI21X1 AOI21X1_502 ( .A(_2739_), .B(_2740_), .C(_2618__bF_buf2), .Y(_2614__21_) );
	NAND2X1 NAND2X1_372 ( .A(_0__22_), .B(_2625__bF_buf1), .Y(_2741_) );
	NAND2X1 NAND2X1_373 ( .A(bounty_synth_22_), .B(_2633__bF_buf1), .Y(_2742_) );
	AOI21X1 AOI21X1_503 ( .A(_2741_), .B(_2742_), .C(_2618__bF_buf1), .Y(_2614__22_) );
	NAND2X1 NAND2X1_374 ( .A(_0__23_), .B(_2625__bF_buf0), .Y(_2743_) );
	NAND2X1 NAND2X1_375 ( .A(bounty_synth_23_), .B(_2633__bF_buf0), .Y(_2744_) );
	AOI21X1 AOI21X1_504 ( .A(_2743_), .B(_2744_), .C(_2618__bF_buf0), .Y(_2614__23_) );
	OAI21X1 OAI21X1_664 ( .A(_2629_), .B(_2630_), .C(RAM_rd_ptr_0_), .Y(_2745_) );
	NAND3X1 NAND3X1_93 ( .A(_2628_), .B(_2623_), .C(_2621_), .Y(_2746_) );
	AOI21X1 AOI21X1_505 ( .A(_2746_), .B(_2745_), .C(_2618__bF_buf6), .Y(_2617__0_) );
	NAND3X1 NAND3X1_94 ( .A(num_entradas[1]), .B(RAM_rd_ptr_0_), .C(comparador_valid_bF_buf0), .Y(_2747_) );
	AOI21X1 AOI21X1_506 ( .A(_2627_), .B(_2747_), .C(_2618__bF_buf5), .Y(_2617__1_) );
	NAND3X1 NAND3X1_95 ( .A(_2623_), .B(_2624_), .C(_2629_), .Y(_2748_) );
	OAI21X1 OAI21X1_665 ( .A(_2629_), .B(_2630_), .C(_1__bF_buf2), .Y(_2749_) );
	AOI21X1 AOI21X1_507 ( .A(_2748_), .B(_2749_), .C(_2618__bF_buf4), .Y(_2615_) );
	DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_bF_buf71), .D(_2615_), .Q(_1_) );
	DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_bF_buf70), .D(_2617__0_), .Q(RAM_rd_ptr_0_) );
	DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_bF_buf69), .D(_2617__1_), .Q(RAM_rd_ptr_1_) );
	DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_bF_buf68), .D(_2614__0_), .Q(_0__0_) );
	DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_bF_buf67), .D(_2614__1_), .Q(_0__1_) );
	DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_bF_buf66), .D(_2614__2_), .Q(_0__2_) );
	DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_bF_buf65), .D(_2614__3_), .Q(_0__3_) );
	DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_bF_buf64), .D(_2614__4_), .Q(_0__4_) );
	DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_bF_buf63), .D(_2614__5_), .Q(_0__5_) );
	DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_bF_buf62), .D(_2614__6_), .Q(_0__6_) );
	DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_bF_buf61), .D(_2614__7_), .Q(_0__7_) );
	DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_bF_buf60), .D(_2614__8_), .Q(_0__8_) );
	DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_bF_buf59), .D(_2614__9_), .Q(_0__9_) );
	DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_bF_buf58), .D(_2614__10_), .Q(_0__10_) );
	DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_bF_buf57), .D(_2614__11_), .Q(_0__11_) );
	DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_bF_buf56), .D(_2614__12_), .Q(_0__12_) );
	DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_bF_buf55), .D(_2614__13_), .Q(_0__13_) );
	DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_bF_buf54), .D(_2614__14_), .Q(_0__14_) );
	DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_bF_buf53), .D(_2614__15_), .Q(_0__15_) );
	DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_bF_buf52), .D(_2614__16_), .Q(_0__16_) );
	DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_bF_buf51), .D(_2614__17_), .Q(_0__17_) );
	DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_bF_buf50), .D(_2614__18_), .Q(_0__18_) );
	DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_bF_buf49), .D(_2614__19_), .Q(_0__19_) );
	DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_bF_buf48), .D(_2614__20_), .Q(_0__20_) );
	DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_bF_buf47), .D(_2614__21_), .Q(_0__21_) );
	DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_bF_buf46), .D(_2614__22_), .Q(_0__22_) );
	DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_bF_buf45), .D(_2614__23_), .Q(_0__23_) );
	DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_bF_buf44), .D(_2616__0_), .Q(_3__0_) );
	DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_bF_buf43), .D(_2616__1_), .Q(_3__1_) );
	DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_bF_buf42), .D(_2616__2_), .Q(_3__2_) );
	DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_bF_buf41), .D(_2616__3_), .Q(_3__3_) );
	DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_bF_buf40), .D(_2616__4_), .Q(_3__4_) );
	DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_bF_buf39), .D(_2616__5_), .Q(_3__5_) );
	DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_bF_buf38), .D(_2616__6_), .Q(_3__6_) );
	DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_bF_buf37), .D(_2616__7_), .Q(_3__7_) );
	DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_bF_buf36), .D(_2616__8_), .Q(_3__8_) );
	DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_bF_buf35), .D(_2616__9_), .Q(_3__9_) );
	DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_bF_buf34), .D(_2616__10_), .Q(_3__10_) );
	DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_bF_buf33), .D(_2616__11_), .Q(_3__11_) );
	DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_bF_buf32), .D(_2616__12_), .Q(_3__12_) );
	DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_bF_buf31), .D(_2616__13_), .Q(_3__13_) );
	DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_bF_buf30), .D(_2616__14_), .Q(_3__14_) );
	DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_bF_buf29), .D(_2616__15_), .Q(_3__15_) );
	DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_bF_buf28), .D(_2616__16_), .Q(_3__16_) );
	DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_bF_buf27), .D(_2616__17_), .Q(_3__17_) );
	DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_bF_buf26), .D(_2616__18_), .Q(_3__18_) );
	DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_bF_buf25), .D(_2616__19_), .Q(_3__19_) );
	DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_bF_buf24), .D(_2616__20_), .Q(_3__20_) );
	DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_bF_buf23), .D(_2616__21_), .Q(_3__21_) );
	DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_bF_buf22), .D(_2616__22_), .Q(_3__22_) );
	DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_bF_buf21), .D(_2616__23_), .Q(_3__23_) );
	DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_bF_buf20), .D(_2616__24_), .Q(_3__24_) );
	DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_bF_buf19), .D(_2616__25_), .Q(_3__25_) );
	DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_bF_buf18), .D(_2616__26_), .Q(_3__26_) );
	DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_bF_buf17), .D(_2616__27_), .Q(_3__27_) );
	DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_bF_buf16), .D(_2616__28_), .Q(_3__28_) );
	DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_bF_buf15), .D(_2616__29_), .Q(_3__29_) );
	DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_bF_buf14), .D(_2616__30_), .Q(_3__30_) );
	DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_bF_buf13), .D(_2616__31_), .Q(_3__31_) );
endmodule
