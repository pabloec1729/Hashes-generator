module hash_synth (target, clk, reset_L, num_entradas, bounty_synth_out, nonce_synth_valido_out, nonce_synth, fin_synth);

input clk;
input reset_L;
output fin_synth;
input [7:0] target;
input [1:0] num_entradas;
output [23:0] bounty_synth_out;
output [31:0] nonce_synth_valido_out;
output [31:0] nonce_synth;

wire vdd = 1'b1;
wire gnd = 1'b0;

	BUFX4 BUFX4_1 ( .A(clk), .Y(clk_hier0_bF_buf9) );
	BUFX4 BUFX4_2 ( .A(clk), .Y(clk_hier0_bF_buf8) );
	BUFX4 BUFX4_3 ( .A(clk), .Y(clk_hier0_bF_buf7) );
	BUFX4 BUFX4_4 ( .A(clk), .Y(clk_hier0_bF_buf6) );
	BUFX4 BUFX4_5 ( .A(clk), .Y(clk_hier0_bF_buf5) );
	BUFX4 BUFX4_6 ( .A(clk), .Y(clk_hier0_bF_buf4) );
	BUFX4 BUFX4_7 ( .A(clk), .Y(clk_hier0_bF_buf3) );
	BUFX4 BUFX4_8 ( .A(clk), .Y(clk_hier0_bF_buf2) );
	BUFX4 BUFX4_9 ( .A(clk), .Y(clk_hier0_bF_buf1) );
	BUFX4 BUFX4_10 ( .A(clk), .Y(clk_hier0_bF_buf0) );
	BUFX2 BUFX2_1 ( .A(reset_L), .Y(reset_L_hier0_bF_buf6) );
	BUFX2 BUFX2_2 ( .A(reset_L), .Y(reset_L_hier0_bF_buf5) );
	BUFX2 BUFX2_3 ( .A(reset_L), .Y(reset_L_hier0_bF_buf4) );
	BUFX2 BUFX2_4 ( .A(reset_L), .Y(reset_L_hier0_bF_buf3) );
	BUFX2 BUFX2_5 ( .A(reset_L), .Y(reset_L_hier0_bF_buf2) );
	BUFX2 BUFX2_6 ( .A(reset_L), .Y(reset_L_hier0_bF_buf1) );
	BUFX2 BUFX2_7 ( .A(reset_L), .Y(reset_L_hier0_bF_buf0) );
	BUFX4 BUFX4_11 ( .A(_92_), .Y(_92__bF_buf6) );
	BUFX2 BUFX2_8 ( .A(_92_), .Y(_92__bF_buf5) );
	BUFX2 BUFX2_9 ( .A(_92_), .Y(_92__bF_buf4) );
	BUFX2 BUFX2_10 ( .A(_92_), .Y(_92__bF_buf3) );
	BUFX2 BUFX2_11 ( .A(_92_), .Y(_92__bF_buf2) );
	BUFX2 BUFX2_12 ( .A(_92_), .Y(_92__bF_buf1) );
	BUFX2 BUFX2_13 ( .A(_92_), .Y(_92__bF_buf0) );
	BUFX2 BUFX2_14 ( .A(_1630_), .Y(_1630__bF_buf4) );
	BUFX2 BUFX2_15 ( .A(_1630_), .Y(_1630__bF_buf3) );
	BUFX2 BUFX2_16 ( .A(_1630_), .Y(_1630__bF_buf2) );
	BUFX2 BUFX2_17 ( .A(_1630_), .Y(_1630__bF_buf1) );
	BUFX2 BUFX2_18 ( .A(_1630_), .Y(_1630__bF_buf0) );
	BUFX4 BUFX4_12 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf113) );
	BUFX4 BUFX4_13 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf112) );
	BUFX4 BUFX4_14 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf111) );
	BUFX4 BUFX4_15 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf110) );
	BUFX4 BUFX4_16 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf109) );
	BUFX4 BUFX4_17 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf108) );
	BUFX4 BUFX4_18 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf107) );
	BUFX4 BUFX4_19 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf106) );
	BUFX4 BUFX4_20 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf105) );
	BUFX4 BUFX4_21 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf104) );
	BUFX4 BUFX4_22 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf103) );
	BUFX4 BUFX4_23 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf102) );
	BUFX4 BUFX4_24 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf101) );
	BUFX4 BUFX4_25 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf100) );
	BUFX4 BUFX4_26 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf99) );
	BUFX4 BUFX4_27 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf98) );
	BUFX4 BUFX4_28 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf97) );
	BUFX4 BUFX4_29 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf96) );
	BUFX4 BUFX4_30 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf95) );
	BUFX4 BUFX4_31 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf94) );
	BUFX4 BUFX4_32 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf93) );
	BUFX4 BUFX4_33 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf92) );
	BUFX4 BUFX4_34 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf91) );
	BUFX4 BUFX4_35 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf90) );
	BUFX4 BUFX4_36 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf89) );
	BUFX4 BUFX4_37 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf88) );
	BUFX4 BUFX4_38 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf87) );
	BUFX4 BUFX4_39 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf86) );
	BUFX4 BUFX4_40 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf85) );
	BUFX4 BUFX4_41 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf84) );
	BUFX4 BUFX4_42 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf83) );
	BUFX4 BUFX4_43 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf82) );
	BUFX4 BUFX4_44 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf81) );
	BUFX4 BUFX4_45 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf80) );
	BUFX4 BUFX4_46 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf79) );
	BUFX4 BUFX4_47 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf78) );
	BUFX4 BUFX4_48 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf77) );
	BUFX4 BUFX4_49 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf76) );
	BUFX4 BUFX4_50 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf75) );
	BUFX4 BUFX4_51 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf74) );
	BUFX4 BUFX4_52 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf73) );
	BUFX4 BUFX4_53 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf72) );
	BUFX4 BUFX4_54 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf71) );
	BUFX4 BUFX4_55 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf70) );
	BUFX4 BUFX4_56 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf69) );
	BUFX4 BUFX4_57 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf68) );
	BUFX4 BUFX4_58 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf67) );
	BUFX4 BUFX4_59 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf66) );
	BUFX4 BUFX4_60 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf65) );
	BUFX4 BUFX4_61 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf64) );
	BUFX4 BUFX4_62 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf63) );
	BUFX4 BUFX4_63 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf62) );
	BUFX4 BUFX4_64 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf61) );
	BUFX4 BUFX4_65 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf60) );
	BUFX4 BUFX4_66 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf59) );
	BUFX4 BUFX4_67 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf58) );
	BUFX4 BUFX4_68 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf57) );
	BUFX4 BUFX4_69 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf56) );
	BUFX4 BUFX4_70 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf55) );
	BUFX4 BUFX4_71 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf54) );
	BUFX4 BUFX4_72 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf53) );
	BUFX4 BUFX4_73 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf52) );
	BUFX4 BUFX4_74 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf51) );
	BUFX4 BUFX4_75 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf50) );
	BUFX4 BUFX4_76 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf49) );
	BUFX4 BUFX4_77 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf48) );
	BUFX4 BUFX4_78 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf47) );
	BUFX4 BUFX4_79 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf46) );
	BUFX4 BUFX4_80 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf45) );
	BUFX4 BUFX4_81 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf44) );
	BUFX4 BUFX4_82 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf43) );
	BUFX4 BUFX4_83 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf42) );
	BUFX4 BUFX4_84 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf41) );
	BUFX4 BUFX4_85 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf40) );
	BUFX4 BUFX4_86 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf39) );
	BUFX4 BUFX4_87 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf38) );
	BUFX4 BUFX4_88 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf37) );
	BUFX4 BUFX4_89 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf36) );
	BUFX4 BUFX4_90 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf35) );
	BUFX4 BUFX4_91 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf34) );
	BUFX4 BUFX4_92 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf33) );
	BUFX4 BUFX4_93 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf32) );
	BUFX4 BUFX4_94 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf31) );
	BUFX4 BUFX4_95 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf30) );
	BUFX4 BUFX4_96 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf29) );
	BUFX4 BUFX4_97 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf28) );
	BUFX4 BUFX4_98 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf27) );
	BUFX4 BUFX4_99 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf26) );
	BUFX4 BUFX4_100 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf25) );
	BUFX4 BUFX4_101 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf24) );
	BUFX4 BUFX4_102 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf23) );
	BUFX4 BUFX4_103 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf22) );
	BUFX4 BUFX4_104 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf21) );
	BUFX4 BUFX4_105 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf20) );
	BUFX4 BUFX4_106 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf19) );
	BUFX4 BUFX4_107 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf18) );
	BUFX4 BUFX4_108 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf17) );
	BUFX4 BUFX4_109 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf16) );
	BUFX4 BUFX4_110 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf15) );
	BUFX4 BUFX4_111 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf14) );
	BUFX4 BUFX4_112 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf13) );
	BUFX4 BUFX4_113 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf12) );
	BUFX4 BUFX4_114 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf11) );
	BUFX4 BUFX4_115 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf10) );
	BUFX4 BUFX4_116 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf9) );
	BUFX4 BUFX4_117 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf8) );
	BUFX4 BUFX4_118 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf7) );
	BUFX4 BUFX4_119 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf6) );
	BUFX4 BUFX4_120 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_121 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_122 ( .A(clk_hier0_bF_buf9), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_123 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_124 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_125 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf0) );
	BUFX2 BUFX2_19 ( .A(_117_), .Y(_117__bF_buf6) );
	BUFX2 BUFX2_20 ( .A(_117_), .Y(_117__bF_buf5) );
	BUFX2 BUFX2_21 ( .A(_117_), .Y(_117__bF_buf4) );
	BUFX2 BUFX2_22 ( .A(_117_), .Y(_117__bF_buf3) );
	BUFX2 BUFX2_23 ( .A(_117_), .Y(_117__bF_buf2) );
	BUFX2 BUFX2_24 ( .A(_117_), .Y(_117__bF_buf1) );
	BUFX2 BUFX2_25 ( .A(_117_), .Y(_117__bF_buf0) );
	BUFX2 BUFX2_26 ( .A(_3022_), .Y(_3022__bF_buf5) );
	BUFX2 BUFX2_27 ( .A(_3022_), .Y(_3022__bF_buf4) );
	BUFX2 BUFX2_28 ( .A(_3022_), .Y(_3022__bF_buf3) );
	BUFX2 BUFX2_29 ( .A(_3022_), .Y(_3022__bF_buf2) );
	BUFX2 BUFX2_30 ( .A(_3022_), .Y(_3022__bF_buf1) );
	BUFX2 BUFX2_31 ( .A(_3022_), .Y(_3022__bF_buf0) );
	BUFX4 BUFX4_126 ( .A(_142_), .Y(_142__bF_buf6) );
	BUFX4 BUFX4_127 ( .A(_142_), .Y(_142__bF_buf5) );
	BUFX4 BUFX4_128 ( .A(_142_), .Y(_142__bF_buf4) );
	BUFX4 BUFX4_129 ( .A(_142_), .Y(_142__bF_buf3) );
	BUFX4 BUFX4_130 ( .A(_142_), .Y(_142__bF_buf2) );
	BUFX4 BUFX4_131 ( .A(_142_), .Y(_142__bF_buf1) );
	BUFX4 BUFX4_132 ( .A(_142_), .Y(_142__bF_buf0) );
	BUFX4 BUFX4_133 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf13) );
	BUFX4 BUFX4_134 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf12) );
	BUFX4 BUFX4_135 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf11) );
	BUFX4 BUFX4_136 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf10) );
	BUFX4 BUFX4_137 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf9) );
	BUFX4 BUFX4_138 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf8) );
	BUFX4 BUFX4_139 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf7) );
	BUFX4 BUFX4_140 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf6) );
	BUFX4 BUFX4_141 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf5) );
	BUFX4 BUFX4_142 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf4) );
	BUFX4 BUFX4_143 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf3) );
	BUFX4 BUFX4_144 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf2) );
	BUFX4 BUFX4_145 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf1) );
	BUFX4 BUFX4_146 ( .A(concatenador_counter_0_), .Y(concatenador_counter_0_bF_buf0) );
	BUFX2 BUFX2_32 ( .A(_3316_), .Y(_3316__bF_buf3) );
	BUFX2 BUFX2_33 ( .A(_3316_), .Y(_3316__bF_buf2) );
	BUFX2 BUFX2_34 ( .A(_3316_), .Y(_3316__bF_buf1) );
	BUFX2 BUFX2_35 ( .A(_3316_), .Y(_3316__bF_buf0) );
	BUFX2 BUFX2_36 ( .A(_3443_), .Y(_3443__bF_buf5) );
	BUFX2 BUFX2_37 ( .A(_3443_), .Y(_3443__bF_buf4) );
	BUFX2 BUFX2_38 ( .A(_3443_), .Y(_3443__bF_buf3) );
	BUFX2 BUFX2_39 ( .A(_3443_), .Y(_3443__bF_buf2) );
	BUFX2 BUFX2_40 ( .A(_3443_), .Y(_3443__bF_buf1) );
	BUFX2 BUFX2_41 ( .A(_3443_), .Y(_3443__bF_buf0) );
	BUFX2 BUFX2_42 ( .A(_5004_), .Y(_5004__bF_buf6) );
	BUFX2 BUFX2_43 ( .A(_5004_), .Y(_5004__bF_buf5) );
	BUFX2 BUFX2_44 ( .A(_5004_), .Y(_5004__bF_buf4) );
	BUFX2 BUFX2_45 ( .A(_5004_), .Y(_5004__bF_buf3) );
	BUFX2 BUFX2_46 ( .A(_5004_), .Y(_5004__bF_buf2) );
	BUFX2 BUFX2_47 ( .A(_5004_), .Y(_5004__bF_buf1) );
	BUFX2 BUFX2_48 ( .A(_5004_), .Y(_5004__bF_buf0) );
	BUFX4 BUFX4_147 ( .A(_4735_), .Y(_4735__bF_buf15) );
	BUFX4 BUFX4_148 ( .A(_4735_), .Y(_4735__bF_buf14) );
	BUFX4 BUFX4_149 ( .A(_4735_), .Y(_4735__bF_buf13) );
	BUFX4 BUFX4_150 ( .A(_4735_), .Y(_4735__bF_buf12) );
	BUFX4 BUFX4_151 ( .A(_4735_), .Y(_4735__bF_buf11) );
	BUFX4 BUFX4_152 ( .A(_4735_), .Y(_4735__bF_buf10) );
	BUFX4 BUFX4_153 ( .A(_4735_), .Y(_4735__bF_buf9) );
	BUFX4 BUFX4_154 ( .A(_4735_), .Y(_4735__bF_buf8) );
	BUFX4 BUFX4_155 ( .A(_4735_), .Y(_4735__bF_buf7) );
	BUFX4 BUFX4_156 ( .A(_4735_), .Y(_4735__bF_buf6) );
	BUFX4 BUFX4_157 ( .A(_4735_), .Y(_4735__bF_buf5) );
	BUFX4 BUFX4_158 ( .A(_4735_), .Y(_4735__bF_buf4) );
	BUFX4 BUFX4_159 ( .A(_4735_), .Y(_4735__bF_buf3) );
	BUFX4 BUFX4_160 ( .A(_4735_), .Y(_4735__bF_buf2) );
	BUFX4 BUFX4_161 ( .A(_4735_), .Y(_4735__bF_buf1) );
	BUFX4 BUFX4_162 ( .A(_4735_), .Y(_4735__bF_buf0) );
	BUFX2 BUFX2_49 ( .A(_4832_), .Y(_4832__bF_buf5) );
	BUFX2 BUFX2_50 ( .A(_4832_), .Y(_4832__bF_buf4) );
	BUFX2 BUFX2_51 ( .A(_4832_), .Y(_4832__bF_buf3) );
	BUFX2 BUFX2_52 ( .A(_4832_), .Y(_4832__bF_buf2) );
	BUFX2 BUFX2_53 ( .A(_4832_), .Y(_4832__bF_buf1) );
	BUFX2 BUFX2_54 ( .A(_4832_), .Y(_4832__bF_buf0) );
	BUFX4 BUFX4_163 ( .A(mux1_sel), .Y(mux1_sel_bF_buf4) );
	BUFX2 BUFX2_55 ( .A(mux1_sel), .Y(mux1_sel_bF_buf3) );
	BUFX2 BUFX2_56 ( .A(mux1_sel), .Y(mux1_sel_bF_buf2) );
	BUFX2 BUFX2_57 ( .A(mux1_sel), .Y(mux1_sel_bF_buf1) );
	BUFX2 BUFX2_58 ( .A(mux1_sel), .Y(mux1_sel_bF_buf0) );
	BUFX2 BUFX2_59 ( .A(RAM_entrada_71_), .Y(RAM_entrada_71_bF_buf3) );
	BUFX2 BUFX2_60 ( .A(RAM_entrada_71_), .Y(RAM_entrada_71_bF_buf2) );
	BUFX2 BUFX2_61 ( .A(RAM_entrada_71_), .Y(RAM_entrada_71_bF_buf1) );
	BUFX2 BUFX2_62 ( .A(RAM_entrada_71_), .Y(RAM_entrada_71_bF_buf0) );
	BUFX2 BUFX2_63 ( .A(_3489_), .Y(_3489__bF_buf3) );
	BUFX2 BUFX2_64 ( .A(_3489_), .Y(_3489__bF_buf2) );
	BUFX2 BUFX2_65 ( .A(_3489_), .Y(_3489__bF_buf1) );
	BUFX2 BUFX2_66 ( .A(_3489_), .Y(_3489__bF_buf0) );
	BUFX2 BUFX2_67 ( .A(_3424_), .Y(_3424__bF_buf3) );
	BUFX2 BUFX2_68 ( .A(_3424_), .Y(_3424__bF_buf2) );
	BUFX2 BUFX2_69 ( .A(_3424_), .Y(_3424__bF_buf1) );
	BUFX2 BUFX2_70 ( .A(_3424_), .Y(_3424__bF_buf0) );
	BUFX2 BUFX2_71 ( .A(_868_), .Y(_868__bF_buf3) );
	BUFX2 BUFX2_72 ( .A(_868_), .Y(_868__bF_buf2) );
	BUFX2 BUFX2_73 ( .A(_868_), .Y(_868__bF_buf1) );
	BUFX2 BUFX2_74 ( .A(_868_), .Y(_868__bF_buf0) );
	BUFX2 BUFX2_75 ( .A(_3442_), .Y(_3442__bF_buf4) );
	BUFX2 BUFX2_76 ( .A(_3442_), .Y(_3442__bF_buf3) );
	BUFX2 BUFX2_77 ( .A(_3442_), .Y(_3442__bF_buf2) );
	BUFX2 BUFX2_78 ( .A(_3442_), .Y(_3442__bF_buf1) );
	BUFX2 BUFX2_79 ( .A(_3442_), .Y(_3442__bF_buf0) );
	BUFX2 BUFX2_80 ( .A(_4269_), .Y(_4269__bF_buf6) );
	BUFX2 BUFX2_81 ( .A(_4269_), .Y(_4269__bF_buf5) );
	BUFX2 BUFX2_82 ( .A(_4269_), .Y(_4269__bF_buf4) );
	BUFX2 BUFX2_83 ( .A(_4269_), .Y(_4269__bF_buf3) );
	BUFX2 BUFX2_84 ( .A(_4269_), .Y(_4269__bF_buf2) );
	BUFX2 BUFX2_85 ( .A(_4269_), .Y(_4269__bF_buf1) );
	BUFX2 BUFX2_86 ( .A(_4269_), .Y(_4269__bF_buf0) );
	BUFX2 BUFX2_87 ( .A(_3333_), .Y(_3333__bF_buf3) );
	BUFX2 BUFX2_88 ( .A(_3333_), .Y(_3333__bF_buf2) );
	BUFX2 BUFX2_89 ( .A(_3333_), .Y(_3333__bF_buf1) );
	BUFX2 BUFX2_90 ( .A(_3333_), .Y(_3333__bF_buf0) );
	BUFX2 BUFX2_91 ( .A(_1506_), .Y(_1506__bF_buf3) );
	BUFX2 BUFX2_92 ( .A(_1506_), .Y(_1506__bF_buf2) );
	BUFX2 BUFX2_93 ( .A(_1506_), .Y(_1506__bF_buf1) );
	BUFX2 BUFX2_94 ( .A(_1506_), .Y(_1506__bF_buf0) );
	BUFX4 BUFX4_164 ( .A(_550_), .Y(_550__bF_buf15) );
	BUFX4 BUFX4_165 ( .A(_550_), .Y(_550__bF_buf14) );
	BUFX4 BUFX4_166 ( .A(_550_), .Y(_550__bF_buf13) );
	BUFX4 BUFX4_167 ( .A(_550_), .Y(_550__bF_buf12) );
	BUFX4 BUFX4_168 ( .A(_550_), .Y(_550__bF_buf11) );
	BUFX4 BUFX4_169 ( .A(_550_), .Y(_550__bF_buf10) );
	BUFX4 BUFX4_170 ( .A(_550_), .Y(_550__bF_buf9) );
	BUFX4 BUFX4_171 ( .A(_550_), .Y(_550__bF_buf8) );
	BUFX4 BUFX4_172 ( .A(_550_), .Y(_550__bF_buf7) );
	BUFX4 BUFX4_173 ( .A(_550_), .Y(_550__bF_buf6) );
	BUFX4 BUFX4_174 ( .A(_550_), .Y(_550__bF_buf5) );
	BUFX4 BUFX4_175 ( .A(_550_), .Y(_550__bF_buf4) );
	BUFX4 BUFX4_176 ( .A(_550_), .Y(_550__bF_buf3) );
	BUFX4 BUFX4_177 ( .A(_550_), .Y(_550__bF_buf2) );
	BUFX4 BUFX4_178 ( .A(_550_), .Y(_550__bF_buf1) );
	BUFX4 BUFX4_179 ( .A(_550_), .Y(_550__bF_buf0) );
	BUFX2 BUFX2_95 ( .A(_1633_), .Y(_1633__bF_buf5) );
	BUFX2 BUFX2_96 ( .A(_1633_), .Y(_1633__bF_buf4) );
	BUFX2 BUFX2_97 ( .A(_1633_), .Y(_1633__bF_buf3) );
	BUFX2 BUFX2_98 ( .A(_1633_), .Y(_1633__bF_buf2) );
	BUFX2 BUFX2_99 ( .A(_1633_), .Y(_1633__bF_buf1) );
	BUFX2 BUFX2_100 ( .A(_1633_), .Y(_1633__bF_buf0) );
	BUFX2 BUFX2_101 ( .A(_53_), .Y(_53__bF_buf6) );
	BUFX2 BUFX2_102 ( .A(_53_), .Y(_53__bF_buf5) );
	BUFX2 BUFX2_103 ( .A(_53_), .Y(_53__bF_buf4) );
	BUFX2 BUFX2_104 ( .A(_53_), .Y(_53__bF_buf3) );
	BUFX2 BUFX2_105 ( .A(_53_), .Y(_53__bF_buf2) );
	BUFX2 BUFX2_106 ( .A(_53_), .Y(_53__bF_buf1) );
	BUFX2 BUFX2_107 ( .A(_53_), .Y(_53__bF_buf0) );
	BUFX2 BUFX2_108 ( .A(concatenador_counter_2d_1_), .Y(concatenador_counter_2d_1_bF_buf6) );
	BUFX2 BUFX2_109 ( .A(concatenador_counter_2d_1_), .Y(concatenador_counter_2d_1_bF_buf5) );
	BUFX4 BUFX4_180 ( .A(concatenador_counter_2d_1_), .Y(concatenador_counter_2d_1_bF_buf4) );
	BUFX2 BUFX2_110 ( .A(concatenador_counter_2d_1_), .Y(concatenador_counter_2d_1_bF_buf3) );
	BUFX2 BUFX2_111 ( .A(concatenador_counter_2d_1_), .Y(concatenador_counter_2d_1_bF_buf2) );
	BUFX2 BUFX2_112 ( .A(concatenador_counter_2d_1_), .Y(concatenador_counter_2d_1_bF_buf1) );
	BUFX2 BUFX2_113 ( .A(concatenador_counter_2d_1_), .Y(concatenador_counter_2d_1_bF_buf0) );
	BUFX2 BUFX2_114 ( .A(comparador_valid), .Y(comparador_valid_bF_buf5) );
	BUFX2 BUFX2_115 ( .A(comparador_valid), .Y(comparador_valid_bF_buf4) );
	BUFX2 BUFX2_116 ( .A(comparador_valid), .Y(comparador_valid_bF_buf3) );
	BUFX2 BUFX2_117 ( .A(comparador_valid), .Y(comparador_valid_bF_buf2) );
	BUFX4 BUFX4_181 ( .A(comparador_valid), .Y(comparador_valid_bF_buf1) );
	BUFX2 BUFX2_118 ( .A(comparador_valid), .Y(comparador_valid_bF_buf0) );
	BUFX2 BUFX2_119 ( .A(_3453_), .Y(_3453__bF_buf3) );
	BUFX2 BUFX2_120 ( .A(_3453_), .Y(_3453__bF_buf2) );
	BUFX2 BUFX2_121 ( .A(_3453_), .Y(_3453__bF_buf1) );
	BUFX2 BUFX2_122 ( .A(_3453_), .Y(_3453__bF_buf0) );
	BUFX4 BUFX4_182 ( .A(_2925_), .Y(_2925__bF_buf15) );
	BUFX4 BUFX4_183 ( .A(_2925_), .Y(_2925__bF_buf14) );
	BUFX4 BUFX4_184 ( .A(_2925_), .Y(_2925__bF_buf13) );
	BUFX4 BUFX4_185 ( .A(_2925_), .Y(_2925__bF_buf12) );
	BUFX4 BUFX4_186 ( .A(_2925_), .Y(_2925__bF_buf11) );
	BUFX4 BUFX4_187 ( .A(_2925_), .Y(_2925__bF_buf10) );
	BUFX4 BUFX4_188 ( .A(_2925_), .Y(_2925__bF_buf9) );
	BUFX4 BUFX4_189 ( .A(_2925_), .Y(_2925__bF_buf8) );
	BUFX4 BUFX4_190 ( .A(_2925_), .Y(_2925__bF_buf7) );
	BUFX4 BUFX4_191 ( .A(_2925_), .Y(_2925__bF_buf6) );
	BUFX4 BUFX4_192 ( .A(_2925_), .Y(_2925__bF_buf5) );
	BUFX4 BUFX4_193 ( .A(_2925_), .Y(_2925__bF_buf4) );
	BUFX4 BUFX4_194 ( .A(_2925_), .Y(_2925__bF_buf3) );
	BUFX4 BUFX4_195 ( .A(_2925_), .Y(_2925__bF_buf2) );
	BUFX4 BUFX4_196 ( .A(_2925_), .Y(_2925__bF_buf1) );
	BUFX4 BUFX4_197 ( .A(_2925_), .Y(_2925__bF_buf0) );
	BUFX2 BUFX2_123 ( .A(_4919_), .Y(_4919__bF_buf4) );
	BUFX2 BUFX2_124 ( .A(_4919_), .Y(_4919__bF_buf3) );
	BUFX2 BUFX2_125 ( .A(_4919_), .Y(_4919__bF_buf2) );
	BUFX2 BUFX2_126 ( .A(_4919_), .Y(_4919__bF_buf1) );
	BUFX2 BUFX2_127 ( .A(_4919_), .Y(_4919__bF_buf0) );
	BUFX2 BUFX2_128 ( .A(_1679_), .Y(_1679__bF_buf3) );
	BUFX2 BUFX2_129 ( .A(_1679_), .Y(_1679__bF_buf2) );
	BUFX2 BUFX2_130 ( .A(_1679_), .Y(_1679__bF_buf1) );
	BUFX2 BUFX2_131 ( .A(_1679_), .Y(_1679__bF_buf0) );
	BUFX4 BUFX4_198 ( .A(_4740_), .Y(_4740__bF_buf13) );
	BUFX4 BUFX4_199 ( .A(_4740_), .Y(_4740__bF_buf12) );
	BUFX4 BUFX4_200 ( .A(_4740_), .Y(_4740__bF_buf11) );
	BUFX4 BUFX4_201 ( .A(_4740_), .Y(_4740__bF_buf10) );
	BUFX4 BUFX4_202 ( .A(_4740_), .Y(_4740__bF_buf9) );
	BUFX4 BUFX4_203 ( .A(_4740_), .Y(_4740__bF_buf8) );
	BUFX4 BUFX4_204 ( .A(_4740_), .Y(_4740__bF_buf7) );
	BUFX4 BUFX4_205 ( .A(_4740_), .Y(_4740__bF_buf6) );
	BUFX4 BUFX4_206 ( .A(_4740_), .Y(_4740__bF_buf5) );
	BUFX4 BUFX4_207 ( .A(_4740_), .Y(_4740__bF_buf4) );
	BUFX4 BUFX4_208 ( .A(_4740_), .Y(_4740__bF_buf3) );
	BUFX4 BUFX4_209 ( .A(_4740_), .Y(_4740__bF_buf2) );
	BUFX4 BUFX4_210 ( .A(_4740_), .Y(_4740__bF_buf1) );
	BUFX4 BUFX4_211 ( .A(_4740_), .Y(_4740__bF_buf0) );
	BUFX4 BUFX4_212 ( .A(_290_), .Y(_290__bF_buf15) );
	BUFX4 BUFX4_213 ( .A(_290_), .Y(_290__bF_buf14) );
	BUFX4 BUFX4_214 ( .A(_290_), .Y(_290__bF_buf13) );
	BUFX4 BUFX4_215 ( .A(_290_), .Y(_290__bF_buf12) );
	BUFX4 BUFX4_216 ( .A(_290_), .Y(_290__bF_buf11) );
	BUFX4 BUFX4_217 ( .A(_290_), .Y(_290__bF_buf10) );
	BUFX4 BUFX4_218 ( .A(_290_), .Y(_290__bF_buf9) );
	BUFX4 BUFX4_219 ( .A(_290_), .Y(_290__bF_buf8) );
	BUFX4 BUFX4_220 ( .A(_290_), .Y(_290__bF_buf7) );
	BUFX4 BUFX4_221 ( .A(_290_), .Y(_290__bF_buf6) );
	BUFX4 BUFX4_222 ( .A(_290_), .Y(_290__bF_buf5) );
	BUFX4 BUFX4_223 ( .A(_290_), .Y(_290__bF_buf4) );
	BUFX4 BUFX4_224 ( .A(_290_), .Y(_290__bF_buf3) );
	BUFX4 BUFX4_225 ( .A(_290_), .Y(_290__bF_buf2) );
	BUFX4 BUFX4_226 ( .A(_290_), .Y(_290__bF_buf1) );
	BUFX4 BUFX4_227 ( .A(_290_), .Y(_290__bF_buf0) );
	BUFX2 BUFX2_132 ( .A(_1614_), .Y(_1614__bF_buf3) );
	BUFX2 BUFX2_133 ( .A(_1614_), .Y(_1614__bF_buf2) );
	BUFX2 BUFX2_134 ( .A(_1614_), .Y(_1614__bF_buf1) );
	BUFX2 BUFX2_135 ( .A(_1614_), .Y(_1614__bF_buf0) );
	BUFX2 BUFX2_136 ( .A(_3439_), .Y(_3439__bF_buf3) );
	BUFX2 BUFX2_137 ( .A(_3439_), .Y(_3439__bF_buf2) );
	BUFX2 BUFX2_138 ( .A(_3439_), .Y(_3439__bF_buf1) );
	BUFX2 BUFX2_139 ( .A(_3439_), .Y(_3439__bF_buf0) );
	BUFX2 BUFX2_140 ( .A(_4997_), .Y(_4997__bF_buf6) );
	BUFX2 BUFX2_141 ( .A(_4997_), .Y(_4997__bF_buf5) );
	BUFX2 BUFX2_142 ( .A(_4997_), .Y(_4997__bF_buf4) );
	BUFX2 BUFX2_143 ( .A(_4997_), .Y(_4997__bF_buf3) );
	BUFX2 BUFX2_144 ( .A(_4997_), .Y(_4997__bF_buf2) );
	BUFX2 BUFX2_145 ( .A(_4997_), .Y(_4997__bF_buf1) );
	BUFX2 BUFX2_146 ( .A(_4997_), .Y(_4997__bF_buf0) );
	BUFX4 BUFX4_228 ( .A(_4733_), .Y(_4733__bF_buf7) );
	BUFX4 BUFX4_229 ( .A(_4733_), .Y(_4733__bF_buf6) );
	BUFX4 BUFX4_230 ( .A(_4733_), .Y(_4733__bF_buf5) );
	BUFX4 BUFX4_231 ( .A(_4733_), .Y(_4733__bF_buf4) );
	BUFX2 BUFX2_147 ( .A(_4733_), .Y(_4733__bF_buf3) );
	BUFX4 BUFX4_232 ( .A(_4733_), .Y(_4733__bF_buf2) );
	BUFX4 BUFX4_233 ( .A(_4733_), .Y(_4733__bF_buf1) );
	BUFX2 BUFX2_148 ( .A(_4733_), .Y(_4733__bF_buf0) );
	BUFX2 BUFX2_149 ( .A(_855_), .Y(_855__bF_buf4) );
	BUFX2 BUFX2_150 ( .A(_855_), .Y(_855__bF_buf3) );
	BUFX2 BUFX2_151 ( .A(_855_), .Y(_855__bF_buf2) );
	BUFX2 BUFX2_152 ( .A(_855_), .Y(_855__bF_buf1) );
	BUFX2 BUFX2_153 ( .A(_855_), .Y(_855__bF_buf0) );
	BUFX2 BUFX2_154 ( .A(_3332_), .Y(_3332__bF_buf3) );
	BUFX2 BUFX2_155 ( .A(_3332_), .Y(_3332__bF_buf2) );
	BUFX2 BUFX2_156 ( .A(_3332_), .Y(_3332__bF_buf1) );
	BUFX2 BUFX2_157 ( .A(_3332_), .Y(_3332__bF_buf0) );
	BUFX2 BUFX2_158 ( .A(_1632_), .Y(_1632__bF_buf4) );
	BUFX2 BUFX2_159 ( .A(_1632_), .Y(_1632__bF_buf3) );
	BUFX2 BUFX2_160 ( .A(_1632_), .Y(_1632__bF_buf2) );
	BUFX2 BUFX2_161 ( .A(_1632_), .Y(_1632__bF_buf1) );
	BUFX2 BUFX2_162 ( .A(_1632_), .Y(_1632__bF_buf0) );
	BUFX2 BUFX2_163 ( .A(mux0_sel), .Y(mux0_sel_bF_buf5) );
	BUFX2 BUFX2_164 ( .A(mux0_sel), .Y(mux0_sel_bF_buf4) );
	BUFX2 BUFX2_165 ( .A(mux0_sel), .Y(mux0_sel_bF_buf3) );
	BUFX2 BUFX2_166 ( .A(mux0_sel), .Y(mux0_sel_bF_buf2) );
	BUFX2 BUFX2_167 ( .A(mux0_sel), .Y(mux0_sel_bF_buf1) );
	BUFX2 BUFX2_168 ( .A(mux0_sel), .Y(mux0_sel_bF_buf0) );
	BUFX4 BUFX4_234 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf12) );
	BUFX4 BUFX4_235 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf11) );
	BUFX4 BUFX4_236 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf10) );
	BUFX4 BUFX4_237 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf9) );
	BUFX4 BUFX4_238 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf8) );
	BUFX4 BUFX4_239 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf7) );
	BUFX4 BUFX4_240 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf6) );
	BUFX4 BUFX4_241 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf5) );
	BUFX4 BUFX4_242 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf4) );
	BUFX4 BUFX4_243 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf3) );
	BUFX4 BUFX4_244 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf2) );
	BUFX4 BUFX4_245 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf1) );
	BUFX4 BUFX4_246 ( .A(concatenador_counter_2d_0_), .Y(concatenador_counter_2d_0_bF_buf0) );
	BUFX2 BUFX2_169 ( .A(_2459_), .Y(_2459__bF_buf6) );
	BUFX2 BUFX2_170 ( .A(_2459_), .Y(_2459__bF_buf5) );
	BUFX2 BUFX2_171 ( .A(_2459_), .Y(_2459__bF_buf4) );
	BUFX2 BUFX2_172 ( .A(_2459_), .Y(_2459__bF_buf3) );
	BUFX2 BUFX2_173 ( .A(_2459_), .Y(_2459__bF_buf2) );
	BUFX2 BUFX2_174 ( .A(_2459_), .Y(_2459__bF_buf1) );
	BUFX2 BUFX2_175 ( .A(_2459_), .Y(_2459__bF_buf0) );
	BUFX2 BUFX2_176 ( .A(_1523_), .Y(_1523__bF_buf3) );
	BUFX2 BUFX2_177 ( .A(_1523_), .Y(_1523__bF_buf2) );
	BUFX2 BUFX2_178 ( .A(_1523_), .Y(_1523__bF_buf1) );
	BUFX2 BUFX2_179 ( .A(_1523_), .Y(_1523__bF_buf0) );
	BUFX2 BUFX2_180 ( .A(_10_), .Y(_10__bF_buf6) );
	BUFX2 BUFX2_181 ( .A(_10_), .Y(_10__bF_buf5) );
	BUFX2 BUFX2_182 ( .A(_10_), .Y(_10__bF_buf4) );
	BUFX2 BUFX2_183 ( .A(_10_), .Y(_10__bF_buf3) );
	BUFX2 BUFX2_184 ( .A(_10_), .Y(_10__bF_buf2) );
	BUFX2 BUFX2_185 ( .A(_10_), .Y(_10__bF_buf1) );
	BUFX2 BUFX2_186 ( .A(_10_), .Y(_10__bF_buf0) );
	BUFX2 BUFX2_187 ( .A(_1_), .Y(_1__bF_buf5) );
	BUFX2 BUFX2_188 ( .A(_1_), .Y(_1__bF_buf4) );
	BUFX2 BUFX2_189 ( .A(_1_), .Y(_1__bF_buf3) );
	BUFX2 BUFX2_190 ( .A(_1_), .Y(_1__bF_buf2) );
	BUFX2 BUFX2_191 ( .A(_1_), .Y(_1__bF_buf1) );
	BUFX2 BUFX2_192 ( .A(_1_), .Y(_1__bF_buf0) );
	BUFX2 BUFX2_193 ( .A(_3440_), .Y(_3440__bF_buf4) );
	BUFX2 BUFX2_194 ( .A(_3440_), .Y(_3440__bF_buf3) );
	BUFX2 BUFX2_195 ( .A(_3440_), .Y(_3440__bF_buf2) );
	BUFX2 BUFX2_196 ( .A(_3440_), .Y(_3440__bF_buf1) );
	BUFX2 BUFX2_197 ( .A(_3440_), .Y(_3440__bF_buf0) );
	BUFX2 BUFX2_198 ( .A(_1643_), .Y(_1643__bF_buf3) );
	BUFX2 BUFX2_199 ( .A(_1643_), .Y(_1643__bF_buf2) );
	BUFX2 BUFX2_200 ( .A(_1643_), .Y(_1643__bF_buf1) );
	BUFX2 BUFX2_201 ( .A(_1643_), .Y(_1643__bF_buf0) );
	BUFX2 BUFX2_202 ( .A(reset_L_hier0_bF_buf6), .Y(reset_L_bF_buf49) );
	BUFX4 BUFX4_247 ( .A(reset_L_hier0_bF_buf5), .Y(reset_L_bF_buf48) );
	BUFX2 BUFX2_203 ( .A(reset_L_hier0_bF_buf4), .Y(reset_L_bF_buf47) );
	BUFX2 BUFX2_204 ( .A(reset_L_hier0_bF_buf3), .Y(reset_L_bF_buf46) );
	BUFX2 BUFX2_205 ( .A(reset_L_hier0_bF_buf2), .Y(reset_L_bF_buf45) );
	BUFX4 BUFX4_248 ( .A(reset_L_hier0_bF_buf1), .Y(reset_L_bF_buf44) );
	BUFX2 BUFX2_206 ( .A(reset_L_hier0_bF_buf0), .Y(reset_L_bF_buf43) );
	BUFX2 BUFX2_207 ( .A(reset_L_hier0_bF_buf6), .Y(reset_L_bF_buf42) );
	BUFX2 BUFX2_208 ( .A(reset_L_hier0_bF_buf5), .Y(reset_L_bF_buf41) );
	BUFX2 BUFX2_209 ( .A(reset_L_hier0_bF_buf4), .Y(reset_L_bF_buf40) );
	BUFX2 BUFX2_210 ( .A(reset_L_hier0_bF_buf3), .Y(reset_L_bF_buf39) );
	BUFX2 BUFX2_211 ( .A(reset_L_hier0_bF_buf2), .Y(reset_L_bF_buf38) );
	BUFX2 BUFX2_212 ( .A(reset_L_hier0_bF_buf1), .Y(reset_L_bF_buf37) );
	BUFX2 BUFX2_213 ( .A(reset_L_hier0_bF_buf0), .Y(reset_L_bF_buf36) );
	BUFX2 BUFX2_214 ( .A(reset_L_hier0_bF_buf6), .Y(reset_L_bF_buf35) );
	BUFX2 BUFX2_215 ( .A(reset_L_hier0_bF_buf5), .Y(reset_L_bF_buf34) );
	BUFX2 BUFX2_216 ( .A(reset_L_hier0_bF_buf4), .Y(reset_L_bF_buf33) );
	BUFX2 BUFX2_217 ( .A(reset_L_hier0_bF_buf3), .Y(reset_L_bF_buf32) );
	BUFX2 BUFX2_218 ( .A(reset_L_hier0_bF_buf2), .Y(reset_L_bF_buf31) );
	BUFX2 BUFX2_219 ( .A(reset_L_hier0_bF_buf1), .Y(reset_L_bF_buf30) );
	BUFX2 BUFX2_220 ( .A(reset_L_hier0_bF_buf0), .Y(reset_L_bF_buf29) );
	BUFX2 BUFX2_221 ( .A(reset_L_hier0_bF_buf6), .Y(reset_L_bF_buf28) );
	BUFX2 BUFX2_222 ( .A(reset_L_hier0_bF_buf5), .Y(reset_L_bF_buf27) );
	BUFX2 BUFX2_223 ( .A(reset_L_hier0_bF_buf4), .Y(reset_L_bF_buf26) );
	BUFX2 BUFX2_224 ( .A(reset_L_hier0_bF_buf3), .Y(reset_L_bF_buf25) );
	BUFX2 BUFX2_225 ( .A(reset_L_hier0_bF_buf2), .Y(reset_L_bF_buf24) );
	BUFX2 BUFX2_226 ( .A(reset_L_hier0_bF_buf1), .Y(reset_L_bF_buf23) );
	BUFX2 BUFX2_227 ( .A(reset_L_hier0_bF_buf0), .Y(reset_L_bF_buf22) );
	BUFX2 BUFX2_228 ( .A(reset_L_hier0_bF_buf6), .Y(reset_L_bF_buf21) );
	BUFX2 BUFX2_229 ( .A(reset_L_hier0_bF_buf5), .Y(reset_L_bF_buf20) );
	BUFX2 BUFX2_230 ( .A(reset_L_hier0_bF_buf4), .Y(reset_L_bF_buf19) );
	BUFX2 BUFX2_231 ( .A(reset_L_hier0_bF_buf3), .Y(reset_L_bF_buf18) );
	BUFX2 BUFX2_232 ( .A(reset_L_hier0_bF_buf2), .Y(reset_L_bF_buf17) );
	BUFX2 BUFX2_233 ( .A(reset_L_hier0_bF_buf1), .Y(reset_L_bF_buf16) );
	BUFX2 BUFX2_234 ( .A(reset_L_hier0_bF_buf0), .Y(reset_L_bF_buf15) );
	BUFX2 BUFX2_235 ( .A(reset_L_hier0_bF_buf6), .Y(reset_L_bF_buf14) );
	BUFX2 BUFX2_236 ( .A(reset_L_hier0_bF_buf5), .Y(reset_L_bF_buf13) );
	BUFX2 BUFX2_237 ( .A(reset_L_hier0_bF_buf4), .Y(reset_L_bF_buf12) );
	BUFX2 BUFX2_238 ( .A(reset_L_hier0_bF_buf3), .Y(reset_L_bF_buf11) );
	BUFX2 BUFX2_239 ( .A(reset_L_hier0_bF_buf2), .Y(reset_L_bF_buf10) );
	BUFX2 BUFX2_240 ( .A(reset_L_hier0_bF_buf1), .Y(reset_L_bF_buf9) );
	BUFX2 BUFX2_241 ( .A(reset_L_hier0_bF_buf0), .Y(reset_L_bF_buf8) );
	BUFX2 BUFX2_242 ( .A(reset_L_hier0_bF_buf6), .Y(reset_L_bF_buf7) );
	BUFX2 BUFX2_243 ( .A(reset_L_hier0_bF_buf5), .Y(reset_L_bF_buf6) );
	BUFX2 BUFX2_244 ( .A(reset_L_hier0_bF_buf4), .Y(reset_L_bF_buf5) );
	BUFX4 BUFX4_249 ( .A(reset_L_hier0_bF_buf3), .Y(reset_L_bF_buf4) );
	BUFX2 BUFX2_245 ( .A(reset_L_hier0_bF_buf2), .Y(reset_L_bF_buf3) );
	BUFX2 BUFX2_246 ( .A(reset_L_hier0_bF_buf1), .Y(reset_L_bF_buf2) );
	BUFX2 BUFX2_247 ( .A(reset_L_hier0_bF_buf0), .Y(reset_L_bF_buf1) );
	BUFX4 BUFX4_250 ( .A(reset_L_hier0_bF_buf6), .Y(reset_L_bF_buf0) );
	BUFX4 BUFX4_251 ( .A(_2930_), .Y(_2930__bF_buf13) );
	BUFX4 BUFX4_252 ( .A(_2930_), .Y(_2930__bF_buf12) );
	BUFX4 BUFX4_253 ( .A(_2930_), .Y(_2930__bF_buf11) );
	BUFX4 BUFX4_254 ( .A(_2930_), .Y(_2930__bF_buf10) );
	BUFX4 BUFX4_255 ( .A(_2930_), .Y(_2930__bF_buf9) );
	BUFX4 BUFX4_256 ( .A(_2930_), .Y(_2930__bF_buf8) );
	BUFX4 BUFX4_257 ( .A(_2930_), .Y(_2930__bF_buf7) );
	BUFX4 BUFX4_258 ( .A(_2930_), .Y(_2930__bF_buf6) );
	BUFX4 BUFX4_259 ( .A(_2930_), .Y(_2930__bF_buf5) );
	BUFX4 BUFX4_260 ( .A(_2930_), .Y(_2930__bF_buf4) );
	BUFX4 BUFX4_261 ( .A(_2930_), .Y(_2930__bF_buf3) );
	BUFX4 BUFX4_262 ( .A(_2930_), .Y(_2930__bF_buf2) );
	BUFX4 BUFX4_263 ( .A(_2930_), .Y(_2930__bF_buf1) );
	BUFX4 BUFX4_264 ( .A(_2930_), .Y(_2930__bF_buf0) );
	BUFX2 BUFX2_248 ( .A(_1629_), .Y(_1629__bF_buf3) );
	BUFX2 BUFX2_249 ( .A(_1629_), .Y(_1629__bF_buf2) );
	BUFX2 BUFX2_250 ( .A(_1629_), .Y(_1629__bF_buf1) );
	BUFX2 BUFX2_251 ( .A(_1629_), .Y(_1629__bF_buf0) );
	BUFX2 BUFX2_252 ( .A(_2923_), .Y(_2923__bF_buf7) );
	BUFX4 BUFX4_265 ( .A(_2923_), .Y(_2923__bF_buf6) );
	BUFX4 BUFX4_266 ( .A(_2923_), .Y(_2923__bF_buf5) );
	BUFX4 BUFX4_267 ( .A(_2923_), .Y(_2923__bF_buf4) );
	BUFX2 BUFX2_253 ( .A(_2923_), .Y(_2923__bF_buf3) );
	BUFX4 BUFX4_268 ( .A(_2923_), .Y(_2923__bF_buf2) );
	BUFX2 BUFX2_254 ( .A(_2923_), .Y(_2923__bF_buf1) );
	BUFX2 BUFX2_255 ( .A(_2923_), .Y(_2923__bF_buf0) );
	BUFX2 BUFX2_256 ( .A(_1522_), .Y(_1522__bF_buf3) );
	BUFX2 BUFX2_257 ( .A(_1522_), .Y(_1522__bF_buf2) );
	BUFX2 BUFX2_258 ( .A(_1522_), .Y(_1522__bF_buf1) );
	BUFX2 BUFX2_259 ( .A(_1522_), .Y(_1522__bF_buf0) );
	BUFX2 BUFX2_260 ( .A(_5012_), .Y(_5012__bF_buf6) );
	BUFX2 BUFX2_261 ( .A(_5012_), .Y(_5012__bF_buf5) );
	BUFX2 BUFX2_262 ( .A(_5012_), .Y(_5012__bF_buf4) );
	BUFX2 BUFX2_263 ( .A(_5012_), .Y(_5012__bF_buf3) );
	BUFX2 BUFX2_264 ( .A(_5012_), .Y(_5012__bF_buf2) );
	BUFX2 BUFX2_265 ( .A(_5012_), .Y(_5012__bF_buf1) );
	BUFX2 BUFX2_266 ( .A(_5012_), .Y(_5012__bF_buf0) );
	BUFX2 BUFX2_267 ( .A(concatenador_counter_1_), .Y(concatenador_counter_1_bF_buf7) );
	BUFX2 BUFX2_268 ( .A(concatenador_counter_1_), .Y(concatenador_counter_1_bF_buf6) );
	BUFX2 BUFX2_269 ( .A(concatenador_counter_1_), .Y(concatenador_counter_1_bF_buf5) );
	BUFX2 BUFX2_270 ( .A(concatenador_counter_1_), .Y(concatenador_counter_1_bF_buf4) );
	BUFX2 BUFX2_271 ( .A(concatenador_counter_1_), .Y(concatenador_counter_1_bF_buf3) );
	BUFX2 BUFX2_272 ( .A(concatenador_counter_1_), .Y(concatenador_counter_1_bF_buf2) );
	BUFX2 BUFX2_273 ( .A(concatenador_counter_1_), .Y(concatenador_counter_1_bF_buf1) );
	BUFX2 BUFX2_274 ( .A(concatenador_counter_1_), .Y(concatenador_counter_1_bF_buf0) );
	BUFX2 BUFX2_275 ( .A(RAM_entrada_84_), .Y(RAM_entrada_84_bF_buf3) );
	BUFX2 BUFX2_276 ( .A(RAM_entrada_84_), .Y(RAM_entrada_84_bF_buf2) );
	BUFX2 BUFX2_277 ( .A(RAM_entrada_84_), .Y(RAM_entrada_84_bF_buf1) );
	BUFX2 BUFX2_278 ( .A(RAM_entrada_84_), .Y(RAM_entrada_84_bF_buf0) );
	OAI22X1 OAI22X1_1 ( .A(_3582_), .B(concatenador_counter_2d_1_bF_buf6), .C(_3580_), .D(_3581_), .Y(_3583_) );
	NAND2X1 NAND2X1_1 ( .A(_3443__bF_buf5), .B(_3583_), .Y(_3584_) );
	AOI21X1 AOI21X1_1 ( .A(_3442__bF_buf4), .B(_3538_), .C(_3453__bF_buf3), .Y(_3585_) );
	NAND3X1 NAND3X1_1 ( .A(_3536_), .B(_3585_), .C(_3584_), .Y(_3586_) );
	NAND3X1 NAND3X1_2 ( .A(_3460_), .B(_3579_), .C(_3586_), .Y(_3587_) );
	NAND2X1 NAND2X1_2 ( .A(_3443__bF_buf4), .B(_3545_), .Y(_3588_) );
	AOI21X1 AOI21X1_2 ( .A(_3440__bF_buf4), .B(_3551_), .C(_3453__bF_buf2), .Y(_3589_) );
	NAND3X1 NAND3X1_3 ( .A(_3549_), .B(_3589_), .C(_3588_), .Y(_3590_) );
	NOR2X1 NOR2X1_1 ( .A(micro_hash_synth_2_W_5__1_), .B(_4733__bF_buf7), .Y(_3591_) );
	OAI21X1 OAI21X1_1 ( .A(concatenador_counter_2d_0_bF_buf12), .B(micro_hash_synth_2_W_4__1_), .C(concatenador_counter_2d_1_bF_buf5), .Y(_3592_) );
	MUX2X1 MUX2X1_1 ( .A(micro_hash_synth_2_W_7__1_), .B(micro_hash_synth_2_W_6__1_), .S(concatenador_counter_2d_0_bF_buf11), .Y(_3593_) );
	OAI22X1 OAI22X1_2 ( .A(_3593_), .B(concatenador_counter_2d_1_bF_buf4), .C(_3591_), .D(_3592_), .Y(_3594_) );
	NAND2X1 NAND2X1_3 ( .A(_3443__bF_buf3), .B(_3594_), .Y(_3595_) );
	AOI21X1 AOI21X1_3 ( .A(_3442__bF_buf3), .B(_3568_), .C(_3489__bF_buf3), .Y(_3596_) );
	NAND3X1 NAND3X1_4 ( .A(_3566_), .B(_3596_), .C(_3595_), .Y(_3597_) );
	NAND3X1 NAND3X1_5 ( .A(_3490_), .B(_3590_), .C(_3597_), .Y(_3598_) );
	INVX1 INVX1_1 ( .A(_3575_), .Y(_3599_) );
	NAND3X1 NAND3X1_6 ( .A(_3599_), .B(_3587_), .C(_3598_), .Y(_3600_) );
	NAND3X1 NAND3X1_7 ( .A(_3576_), .B(_3600_), .C(_3508_), .Y(_3601_) );
	INVX1 INVX1_2 ( .A(_3601_), .Y(_3602_) );
	INVX2 INVX2_1 ( .A(_3505_), .Y(_3603_) );
	NAND2X1 NAND2X1_4 ( .A(_3600_), .B(_3576_), .Y(_3604_) );
	INVX1 INVX1_3 ( .A(_3604_), .Y(_3605_) );
	OAI21X1 OAI21X1_2 ( .A(_3605_), .B(_3508_), .C(_3603_), .Y(_3606_) );
	AOI21X1 AOI21X1_4 ( .A(micro_hash_synth_2_c_1_), .B(_3436_), .C(_3332__bF_buf3), .Y(_3607_) );
	OAI21X1 OAI21X1_3 ( .A(_3606_), .B(_3602_), .C(_3607_), .Y(_3050__1_) );
	AOI21X1 AOI21X1_5 ( .A(_3587_), .B(_3598_), .C(_3599_), .Y(_3608_) );
	NOR2X1 NOR2X1_2 ( .A(micro_hash_synth_2_W_21__2_), .B(_4733__bF_buf6), .Y(_3609_) );
	OAI21X1 OAI21X1_4 ( .A(concatenador_counter_2d_0_bF_buf10), .B(micro_hash_synth_2_W_20__2_), .C(concatenador_counter_2d_1_bF_buf3), .Y(_3610_) );
	MUX2X1 MUX2X1_2 ( .A(micro_hash_synth_2_W_23__2_), .B(micro_hash_synth_2_W_22__2_), .S(concatenador_counter_2d_0_bF_buf9), .Y(_3611_) );
	OAI22X1 OAI22X1_3 ( .A(_3611_), .B(concatenador_counter_2d_1_bF_buf2), .C(_3609_), .D(_3610_), .Y(_3612_) );
	NAND2X1 NAND2X1_5 ( .A(_3443__bF_buf2), .B(_3612_), .Y(_3613_) );
	INVX1 INVX1_4 ( .A(micro_hash_synth_2_W_18__2_), .Y(_3614_) );
	NAND2X1 NAND2X1_6 ( .A(concatenador_counter_2d_0_bF_buf8), .B(micro_hash_synth_2_W_19__2_), .Y(_3615_) );
	OAI21X1 OAI21X1_5 ( .A(_3614_), .B(concatenador_counter_2d_0_bF_buf7), .C(_3615_), .Y(_3616_) );
	NAND2X1 NAND2X1_7 ( .A(_3442__bF_buf2), .B(_3616_), .Y(_3617_) );
	INVX1 INVX1_5 ( .A(micro_hash_synth_2_W_16__2_), .Y(_3618_) );
	NAND2X1 NAND2X1_8 ( .A(concatenador_counter_2d_0_bF_buf6), .B(micro_hash_synth_2_W_17__2_), .Y(_3619_) );
	OAI21X1 OAI21X1_6 ( .A(_3618_), .B(concatenador_counter_2d_0_bF_buf5), .C(_3619_), .Y(_3620_) );
	AOI21X1 AOI21X1_6 ( .A(_3440__bF_buf3), .B(_3620_), .C(_3489__bF_buf2), .Y(_3621_) );
	NAND3X1 NAND3X1_8 ( .A(_3617_), .B(_3621_), .C(_3613_), .Y(_3622_) );
	NOR2X1 NOR2X1_3 ( .A(micro_hash_synth_2_W_29__2_), .B(_4733__bF_buf5), .Y(_3623_) );
	OAI21X1 OAI21X1_7 ( .A(concatenador_counter_2d_0_bF_buf4), .B(micro_hash_synth_2_W_28__2_), .C(concatenador_counter_2d_1_bF_buf1), .Y(_3624_) );
	NOR2X1 NOR2X1_4 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_30__2_), .Y(_3625_) );
	OAI21X1 OAI21X1_8 ( .A(_4733__bF_buf4), .B(micro_hash_synth_2_W_31__2_), .C(_3439__bF_buf3), .Y(_3626_) );
	OAI22X1 OAI22X1_4 ( .A(_3623_), .B(_3624_), .C(_3626_), .D(_3625_), .Y(_3627_) );
	NAND2X1 NAND2X1_9 ( .A(_3443__bF_buf1), .B(_3627_), .Y(_3628_) );
	INVX1 INVX1_6 ( .A(micro_hash_synth_2_W_24__2_), .Y(_3629_) );
	NAND2X1 NAND2X1_10 ( .A(concatenador_counter_2d_0_bF_buf2), .B(micro_hash_synth_2_W_25__2_), .Y(_3630_) );
	OAI21X1 OAI21X1_9 ( .A(_3629_), .B(concatenador_counter_2d_0_bF_buf1), .C(_3630_), .Y(_3631_) );
	NAND2X1 NAND2X1_11 ( .A(_3440__bF_buf2), .B(_3631_), .Y(_3632_) );
	NAND2X1 NAND2X1_12 ( .A(concatenador_counter_2d_0_bF_buf0), .B(micro_hash_synth_2_W_27__2_), .Y(_3633_) );
	OAI21X1 OAI21X1_10 ( .A(_4748_), .B(concatenador_counter_2d_0_bF_buf12), .C(_3633_), .Y(_3634_) );
	AOI21X1 AOI21X1_7 ( .A(_3442__bF_buf1), .B(_3634_), .C(_3453__bF_buf1), .Y(_3635_) );
	NAND3X1 NAND3X1_9 ( .A(_3632_), .B(_3635_), .C(_3628_), .Y(_3636_) );
	NAND3X1 NAND3X1_10 ( .A(_3460_), .B(_3622_), .C(_3636_), .Y(_3637_) );
	NOR2X1 NOR2X1_5 ( .A(micro_hash_synth_2_W_13__2_), .B(_4733__bF_buf3), .Y(_3638_) );
	OAI21X1 OAI21X1_11 ( .A(concatenador_counter_2d_0_bF_buf11), .B(micro_hash_synth_2_W_12__2_), .C(concatenador_counter_2d_1_bF_buf0), .Y(_3639_) );
	MUX2X1 MUX2X1_3 ( .A(micro_hash_synth_2_W_15__2_), .B(micro_hash_synth_2_W_14__2_), .S(concatenador_counter_2d_0_bF_buf10), .Y(_3640_) );
	OAI22X1 OAI22X1_5 ( .A(_3640_), .B(concatenador_counter_2d_1_bF_buf6), .C(_3638_), .D(_3639_), .Y(_3641_) );
	NAND2X1 NAND2X1_13 ( .A(_3443__bF_buf0), .B(_3641_), .Y(_3642_) );
	NAND2X1 NAND2X1_14 ( .A(concatenador_counter_2d_0_bF_buf9), .B(micro_hash_synth_2_W_9__2_), .Y(_3643_) );
	OAI21X1 OAI21X1_12 ( .A(_4804_), .B(concatenador_counter_2d_0_bF_buf8), .C(_3643_), .Y(_3644_) );
	NAND2X1 NAND2X1_15 ( .A(_3440__bF_buf1), .B(_3644_), .Y(_3645_) );
	INVX1 INVX1_7 ( .A(micro_hash_synth_2_W_10__2_), .Y(_3646_) );
	NAND2X1 NAND2X1_16 ( .A(concatenador_counter_2d_0_bF_buf7), .B(micro_hash_synth_2_W_11__2_), .Y(_3647_) );
	OAI21X1 OAI21X1_13 ( .A(_3646_), .B(concatenador_counter_2d_0_bF_buf6), .C(_3647_), .Y(_3648_) );
	AOI21X1 AOI21X1_8 ( .A(_3442__bF_buf0), .B(_3648_), .C(_3453__bF_buf0), .Y(_3649_) );
	NAND3X1 NAND3X1_11 ( .A(_3645_), .B(_3649_), .C(_3642_), .Y(_3650_) );
	NOR2X1 NOR2X1_6 ( .A(micro_hash_synth_2_W_5__2_), .B(_4733__bF_buf2), .Y(_3651_) );
	OAI21X1 OAI21X1_14 ( .A(concatenador_counter_2d_0_bF_buf5), .B(micro_hash_synth_2_W_4__2_), .C(concatenador_counter_2d_1_bF_buf5), .Y(_3652_) );
	NOR2X1 NOR2X1_7 ( .A(concatenador_counter_2d_0_bF_buf4), .B(micro_hash_synth_2_W_6__2_), .Y(_3653_) );
	OAI21X1 OAI21X1_15 ( .A(_4733__bF_buf1), .B(micro_hash_synth_2_W_7__2_), .C(_3439__bF_buf2), .Y(_3654_) );
	OAI22X1 OAI22X1_6 ( .A(_3651_), .B(_3652_), .C(_3654_), .D(_3653_), .Y(_3655_) );
	NAND2X1 NAND2X1_17 ( .A(_3443__bF_buf5), .B(_3655_), .Y(_3656_) );
	NAND2X1 NAND2X1_18 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_1__2_), .Y(_3657_) );
	OAI21X1 OAI21X1_16 ( .A(_4843_), .B(concatenador_counter_2d_0_bF_buf2), .C(_3657_), .Y(_3658_) );
	NAND2X1 NAND2X1_19 ( .A(_3440__bF_buf0), .B(_3658_), .Y(_3659_) );
	NAND2X1 NAND2X1_20 ( .A(concatenador_counter_2d_0_bF_buf1), .B(micro_hash_synth_2_W_3__2_), .Y(_3660_) );
	OAI21X1 OAI21X1_17 ( .A(_4851_), .B(concatenador_counter_2d_0_bF_buf0), .C(_3660_), .Y(_3661_) );
	AOI21X1 AOI21X1_9 ( .A(_3442__bF_buf4), .B(_3661_), .C(_3489__bF_buf1), .Y(_3662_) );
	NAND3X1 NAND3X1_12 ( .A(_3659_), .B(_3662_), .C(_3656_), .Y(_3663_) );
	NAND3X1 NAND3X1_13 ( .A(_3490_), .B(_3650_), .C(_3663_), .Y(_3664_) );
	NAND2X1 NAND2X1_21 ( .A(micro_hash_synth_2_k_2_), .B(micro_hash_synth_2_x_2_), .Y(_3665_) );
	INVX1 INVX1_8 ( .A(micro_hash_synth_2_x_2_), .Y(_3666_) );
	NAND2X1 NAND2X1_22 ( .A(_3428_), .B(_3666_), .Y(_3667_) );
	AND2X2 AND2X2_1 ( .A(_3667_), .B(_3665_), .Y(_3668_) );
	INVX1 INVX1_9 ( .A(_3668_), .Y(_3669_) );
	AOI21X1 AOI21X1_10 ( .A(_3637_), .B(_3664_), .C(_3669_), .Y(_3670_) );
	NAND2X1 NAND2X1_23 ( .A(_3440__bF_buf4), .B(_3620_), .Y(_3671_) );
	NAND3X1 NAND3X1_14 ( .A(_3453__bF_buf3), .B(_3617_), .C(_3671_), .Y(_3672_) );
	AOI21X1 AOI21X1_11 ( .A(_3443__bF_buf4), .B(_3612_), .C(_3672_), .Y(_3673_) );
	INVX1 INVX1_10 ( .A(micro_hash_synth_2_W_29__2_), .Y(_3674_) );
	NAND2X1 NAND2X1_24 ( .A(concatenador_counter_2d_0_bF_buf12), .B(_3674_), .Y(_3675_) );
	OR2X2 OR2X2_1 ( .A(concatenador_counter_2d_0_bF_buf11), .B(micro_hash_synth_2_W_28__2_), .Y(_3676_) );
	NAND3X1 NAND3X1_15 ( .A(concatenador_counter_2d_1_bF_buf4), .B(_3676_), .C(_3675_), .Y(_3677_) );
	OR2X2 OR2X2_2 ( .A(concatenador_counter_2d_0_bF_buf10), .B(micro_hash_synth_2_W_30__2_), .Y(_3678_) );
	INVX1 INVX1_11 ( .A(micro_hash_synth_2_W_31__2_), .Y(_3679_) );
	NAND2X1 NAND2X1_25 ( .A(concatenador_counter_2d_0_bF_buf9), .B(_3679_), .Y(_3680_) );
	NAND3X1 NAND3X1_16 ( .A(_3439__bF_buf1), .B(_3678_), .C(_3680_), .Y(_3681_) );
	AOI21X1 AOI21X1_12 ( .A(_3677_), .B(_3681_), .C(_3523_), .Y(_3682_) );
	NAND2X1 NAND2X1_26 ( .A(_3442__bF_buf3), .B(_3634_), .Y(_3683_) );
	NAND3X1 NAND3X1_17 ( .A(_3489__bF_buf0), .B(_3632_), .C(_3683_), .Y(_3684_) );
	OAI21X1 OAI21X1_18 ( .A(_3684_), .B(_3682_), .C(_3460_), .Y(_3685_) );
	NAND2X1 NAND2X1_27 ( .A(_3442__bF_buf2), .B(_3648_), .Y(_3686_) );
	NAND3X1 NAND3X1_18 ( .A(_3489__bF_buf3), .B(_3645_), .C(_3686_), .Y(_3687_) );
	AOI21X1 AOI21X1_13 ( .A(_3443__bF_buf3), .B(_3641_), .C(_3687_), .Y(_3688_) );
	INVX1 INVX1_12 ( .A(micro_hash_synth_2_W_5__2_), .Y(_3689_) );
	NAND2X1 NAND2X1_28 ( .A(concatenador_counter_2d_0_bF_buf8), .B(_3689_), .Y(_3690_) );
	OR2X2 OR2X2_3 ( .A(concatenador_counter_2d_0_bF_buf7), .B(micro_hash_synth_2_W_4__2_), .Y(_3691_) );
	NAND3X1 NAND3X1_19 ( .A(concatenador_counter_2d_1_bF_buf3), .B(_3691_), .C(_3690_), .Y(_3692_) );
	OR2X2 OR2X2_4 ( .A(concatenador_counter_2d_0_bF_buf6), .B(micro_hash_synth_2_W_6__2_), .Y(_3693_) );
	INVX1 INVX1_13 ( .A(micro_hash_synth_2_W_7__2_), .Y(_3694_) );
	NAND2X1 NAND2X1_29 ( .A(concatenador_counter_2d_0_bF_buf5), .B(_3694_), .Y(_3695_) );
	NAND3X1 NAND3X1_20 ( .A(_3439__bF_buf0), .B(_3693_), .C(_3695_), .Y(_3696_) );
	AOI21X1 AOI21X1_14 ( .A(_3692_), .B(_3696_), .C(_3523_), .Y(_3697_) );
	NAND2X1 NAND2X1_30 ( .A(_3442__bF_buf1), .B(_3661_), .Y(_3698_) );
	NAND3X1 NAND3X1_21 ( .A(_3453__bF_buf2), .B(_3659_), .C(_3698_), .Y(_3699_) );
	OAI21X1 OAI21X1_19 ( .A(_3699_), .B(_3697_), .C(_3490_), .Y(_3700_) );
	OAI22X1 OAI22X1_7 ( .A(_3685_), .B(_3673_), .C(_3688_), .D(_3700_), .Y(_3701_) );
	NOR2X1 NOR2X1_8 ( .A(_3668_), .B(_3701_), .Y(_3702_) );
	OAI22X1 OAI22X1_8 ( .A(_3573_), .B(_3608_), .C(_3702_), .D(_3670_), .Y(_3703_) );
	AOI21X1 AOI21X1_15 ( .A(_3575_), .B(_3572_), .C(_3573_), .Y(_3704_) );
	NAND2X1 NAND2X1_31 ( .A(_3668_), .B(_3701_), .Y(_3705_) );
	NAND3X1 NAND3X1_22 ( .A(_3669_), .B(_3637_), .C(_3664_), .Y(_3706_) );
	NAND3X1 NAND3X1_23 ( .A(_3705_), .B(_3706_), .C(_3704_), .Y(_3707_) );
	NAND2X1 NAND2X1_32 ( .A(_3703_), .B(_3707_), .Y(_3708_) );
	NOR2X1 NOR2X1_9 ( .A(_3602_), .B(_3708_), .Y(_3709_) );
	AOI21X1 AOI21X1_16 ( .A(_3703_), .B(_3707_), .C(_3601_), .Y(_3710_) );
	INVX1 INVX1_14 ( .A(_3710_), .Y(_3711_) );
	NAND2X1 NAND2X1_33 ( .A(_3603_), .B(_3711_), .Y(_3712_) );
	AOI21X1 AOI21X1_17 ( .A(micro_hash_synth_2_c_2_), .B(_3436_), .C(_3332__bF_buf2), .Y(_3713_) );
	OAI21X1 OAI21X1_20 ( .A(_3712_), .B(_3709_), .C(_3713_), .Y(_3050__2_) );
	NAND2X1 NAND2X1_34 ( .A(_3705_), .B(_3706_), .Y(_3714_) );
	NOR2X1 NOR2X1_10 ( .A(_3704_), .B(_3714_), .Y(_3715_) );
	NOR2X1 NOR2X1_11 ( .A(_3715_), .B(_3710_), .Y(_3716_) );
	AOI21X1 AOI21X1_18 ( .A(micro_hash_synth_2_k_2_), .B(micro_hash_synth_2_x_2_), .C(_3670_), .Y(_3717_) );
	NAND2X1 NAND2X1_35 ( .A(micro_hash_synth_2_k_3_), .B(micro_hash_synth_2_x_3_), .Y(_3718_) );
	INVX1 INVX1_15 ( .A(micro_hash_synth_2_x_3_), .Y(_3719_) );
	NAND2X1 NAND2X1_36 ( .A(_3429_), .B(_3719_), .Y(_3720_) );
	AND2X2 AND2X2_2 ( .A(_3720_), .B(_3718_), .Y(_3721_) );
	INVX1 INVX1_16 ( .A(_3721_), .Y(_3722_) );
	NOR2X1 NOR2X1_12 ( .A(micro_hash_synth_2_W_29__3_), .B(_4733__bF_buf0), .Y(_3723_) );
	OAI21X1 OAI21X1_21 ( .A(concatenador_counter_2d_0_bF_buf4), .B(micro_hash_synth_2_W_28__3_), .C(concatenador_counter_2d_1_bF_buf2), .Y(_3724_) );
	NOR2X1 NOR2X1_13 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_30__3_), .Y(_3725_) );
	OAI21X1 OAI21X1_22 ( .A(_4733__bF_buf7), .B(micro_hash_synth_2_W_31__3_), .C(_3439__bF_buf3), .Y(_3726_) );
	OAI22X1 OAI22X1_9 ( .A(_3723_), .B(_3724_), .C(_3726_), .D(_3725_), .Y(_3727_) );
	NAND2X1 NAND2X1_37 ( .A(_3443__bF_buf2), .B(_3727_), .Y(_3728_) );
	INVX1 INVX1_17 ( .A(micro_hash_synth_2_W_24__3_), .Y(_3729_) );
	NAND2X1 NAND2X1_38 ( .A(concatenador_counter_2d_0_bF_buf2), .B(micro_hash_synth_2_W_25__3_), .Y(_3730_) );
	OAI21X1 OAI21X1_23 ( .A(_3729_), .B(concatenador_counter_2d_0_bF_buf1), .C(_3730_), .Y(_3731_) );
	NAND2X1 NAND2X1_39 ( .A(_3440__bF_buf3), .B(_3731_), .Y(_3732_) );
	NAND2X1 NAND2X1_40 ( .A(concatenador_counter_2d_0_bF_buf0), .B(micro_hash_synth_2_W_27__3_), .Y(_3733_) );
	OAI21X1 OAI21X1_24 ( .A(_4753_), .B(concatenador_counter_2d_0_bF_buf12), .C(_3733_), .Y(_3734_) );
	NAND2X1 NAND2X1_41 ( .A(_3442__bF_buf0), .B(_3734_), .Y(_3735_) );
	AND2X2 AND2X2_3 ( .A(_3732_), .B(_3735_), .Y(_3736_) );
	AOI21X1 AOI21X1_19 ( .A(_3728_), .B(_3736_), .C(_3453__bF_buf1), .Y(_3737_) );
	NOR2X1 NOR2X1_14 ( .A(micro_hash_synth_2_W_21__3_), .B(_4733__bF_buf6), .Y(_3738_) );
	OAI21X1 OAI21X1_25 ( .A(concatenador_counter_2d_0_bF_buf11), .B(micro_hash_synth_2_W_20__3_), .C(concatenador_counter_2d_1_bF_buf1), .Y(_3739_) );
	NOR2X1 NOR2X1_15 ( .A(concatenador_counter_2d_0_bF_buf10), .B(micro_hash_synth_2_W_22__3_), .Y(_3740_) );
	OAI21X1 OAI21X1_26 ( .A(_4733__bF_buf5), .B(micro_hash_synth_2_W_23__3_), .C(_3439__bF_buf2), .Y(_3741_) );
	OAI22X1 OAI22X1_10 ( .A(_3738_), .B(_3739_), .C(_3741_), .D(_3740_), .Y(_3742_) );
	NAND2X1 NAND2X1_42 ( .A(_3443__bF_buf1), .B(_3742_), .Y(_3743_) );
	INVX1 INVX1_18 ( .A(micro_hash_synth_2_W_18__3_), .Y(_3744_) );
	NAND2X1 NAND2X1_43 ( .A(concatenador_counter_2d_0_bF_buf9), .B(micro_hash_synth_2_W_19__3_), .Y(_3745_) );
	OAI21X1 OAI21X1_27 ( .A(_3744_), .B(concatenador_counter_2d_0_bF_buf8), .C(_3745_), .Y(_3746_) );
	NAND2X1 NAND2X1_44 ( .A(_3442__bF_buf4), .B(_3746_), .Y(_3747_) );
	INVX1 INVX1_19 ( .A(micro_hash_synth_2_W_16__3_), .Y(_3748_) );
	NAND2X1 NAND2X1_45 ( .A(concatenador_counter_2d_0_bF_buf7), .B(micro_hash_synth_2_W_17__3_), .Y(_3749_) );
	OAI21X1 OAI21X1_28 ( .A(_3748_), .B(concatenador_counter_2d_0_bF_buf6), .C(_3749_), .Y(_3750_) );
	NAND2X1 NAND2X1_46 ( .A(_3440__bF_buf2), .B(_3750_), .Y(_3751_) );
	AND2X2 AND2X2_4 ( .A(_3747_), .B(_3751_), .Y(_3752_) );
	AOI21X1 AOI21X1_20 ( .A(_3743_), .B(_3752_), .C(_3489__bF_buf2), .Y(_3753_) );
	OAI21X1 OAI21X1_29 ( .A(_3737_), .B(_3753_), .C(_3460_), .Y(_3754_) );
	NOR2X1 NOR2X1_16 ( .A(micro_hash_synth_2_W_13__3_), .B(_4733__bF_buf4), .Y(_3755_) );
	OAI21X1 OAI21X1_30 ( .A(concatenador_counter_2d_0_bF_buf5), .B(micro_hash_synth_2_W_12__3_), .C(concatenador_counter_2d_1_bF_buf0), .Y(_3756_) );
	NOR2X1 NOR2X1_17 ( .A(concatenador_counter_2d_0_bF_buf4), .B(micro_hash_synth_2_W_14__3_), .Y(_3757_) );
	OAI21X1 OAI21X1_31 ( .A(_4733__bF_buf3), .B(micro_hash_synth_2_W_15__3_), .C(_3439__bF_buf1), .Y(_3758_) );
	OAI22X1 OAI22X1_11 ( .A(_3755_), .B(_3756_), .C(_3758_), .D(_3757_), .Y(_3759_) );
	NAND2X1 NAND2X1_47 ( .A(_3443__bF_buf0), .B(_3759_), .Y(_3760_) );
	INVX1 INVX1_20 ( .A(micro_hash_synth_2_W_10__3_), .Y(_3761_) );
	NAND2X1 NAND2X1_48 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_11__3_), .Y(_3762_) );
	OAI21X1 OAI21X1_32 ( .A(_3761_), .B(concatenador_counter_2d_0_bF_buf2), .C(_3762_), .Y(_3763_) );
	NAND2X1 NAND2X1_49 ( .A(_3442__bF_buf3), .B(_3763_), .Y(_3764_) );
	NAND2X1 NAND2X1_50 ( .A(concatenador_counter_2d_0_bF_buf1), .B(micro_hash_synth_2_W_9__3_), .Y(_3765_) );
	OAI21X1 OAI21X1_33 ( .A(_4806_), .B(concatenador_counter_2d_0_bF_buf0), .C(_3765_), .Y(_3766_) );
	AOI21X1 AOI21X1_21 ( .A(_3440__bF_buf1), .B(_3766_), .C(_3453__bF_buf0), .Y(_3767_) );
	NAND3X1 NAND3X1_24 ( .A(_3764_), .B(_3767_), .C(_3760_), .Y(_3768_) );
	NOR2X1 NOR2X1_18 ( .A(micro_hash_synth_2_W_5__3_), .B(_4733__bF_buf2), .Y(_3769_) );
	OAI21X1 OAI21X1_34 ( .A(concatenador_counter_2d_0_bF_buf12), .B(micro_hash_synth_2_W_4__3_), .C(concatenador_counter_2d_1_bF_buf6), .Y(_3770_) );
	MUX2X1 MUX2X1_4 ( .A(micro_hash_synth_2_W_7__3_), .B(micro_hash_synth_2_W_6__3_), .S(concatenador_counter_2d_0_bF_buf11), .Y(_3771_) );
	OAI22X1 OAI22X1_12 ( .A(_3771_), .B(concatenador_counter_2d_1_bF_buf5), .C(_3769_), .D(_3770_), .Y(_3772_) );
	AND2X2 AND2X2_5 ( .A(_3772_), .B(_3443__bF_buf5), .Y(_3773_) );
	NAND2X1 NAND2X1_51 ( .A(concatenador_counter_2d_0_bF_buf10), .B(micro_hash_synth_2_W_1__3_), .Y(_3774_) );
	OAI21X1 OAI21X1_35 ( .A(_4844_), .B(concatenador_counter_2d_0_bF_buf9), .C(_3774_), .Y(_3775_) );
	NAND2X1 NAND2X1_52 ( .A(_3440__bF_buf0), .B(_3775_), .Y(_3776_) );
	NAND2X1 NAND2X1_53 ( .A(concatenador_counter_2d_0_bF_buf8), .B(micro_hash_synth_2_W_3__3_), .Y(_3777_) );
	OAI21X1 OAI21X1_36 ( .A(_4852_), .B(concatenador_counter_2d_0_bF_buf7), .C(_3777_), .Y(_3778_) );
	NAND2X1 NAND2X1_54 ( .A(_3442__bF_buf2), .B(_3778_), .Y(_3779_) );
	NAND3X1 NAND3X1_25 ( .A(_3453__bF_buf3), .B(_3776_), .C(_3779_), .Y(_3780_) );
	OR2X2 OR2X2_5 ( .A(_3773_), .B(_3780_), .Y(_3781_) );
	NAND3X1 NAND3X1_26 ( .A(_3490_), .B(_3768_), .C(_3781_), .Y(_3782_) );
	NAND3X1 NAND3X1_27 ( .A(_3722_), .B(_3754_), .C(_3782_), .Y(_3783_) );
	AND2X2 AND2X2_6 ( .A(_3742_), .B(_3443__bF_buf4), .Y(_3784_) );
	NAND3X1 NAND3X1_28 ( .A(_3453__bF_buf2), .B(_3747_), .C(_3751_), .Y(_3785_) );
	AND2X2 AND2X2_7 ( .A(_3727_), .B(_3443__bF_buf3), .Y(_3786_) );
	NAND3X1 NAND3X1_29 ( .A(_3489__bF_buf1), .B(_3732_), .C(_3735_), .Y(_3787_) );
	OAI22X1 OAI22X1_13 ( .A(_3784_), .B(_3785_), .C(_3786_), .D(_3787_), .Y(_3788_) );
	NAND2X1 NAND2X1_55 ( .A(_3460_), .B(_3788_), .Y(_3789_) );
	AND2X2 AND2X2_8 ( .A(_3759_), .B(_3443__bF_buf2), .Y(_3790_) );
	NAND2X1 NAND2X1_56 ( .A(_3440__bF_buf4), .B(_3766_), .Y(_3791_) );
	NAND3X1 NAND3X1_30 ( .A(_3489__bF_buf0), .B(_3764_), .C(_3791_), .Y(_3792_) );
	OAI22X1 OAI22X1_14 ( .A(_3773_), .B(_3780_), .C(_3790_), .D(_3792_), .Y(_3793_) );
	NAND2X1 NAND2X1_57 ( .A(_3490_), .B(_3793_), .Y(_3794_) );
	NAND3X1 NAND3X1_31 ( .A(_3721_), .B(_3794_), .C(_3789_), .Y(_3795_) );
	NAND2X1 NAND2X1_58 ( .A(_3795_), .B(_3783_), .Y(_3796_) );
	NAND2X1 NAND2X1_59 ( .A(_3717_), .B(_3796_), .Y(_3797_) );
	OR2X2 OR2X2_6 ( .A(_3796_), .B(_3717_), .Y(_3798_) );
	NAND2X1 NAND2X1_60 ( .A(_3797_), .B(_3798_), .Y(_3799_) );
	AOI21X1 AOI21X1_22 ( .A(_3799_), .B(_3716_), .C(_3505_), .Y(_3800_) );
	OAI21X1 OAI21X1_37 ( .A(_3716_), .B(_3799_), .C(_3800_), .Y(_3801_) );
	AOI21X1 AOI21X1_23 ( .A(micro_hash_synth_2_c_3_), .B(_3436_), .C(_3332__bF_buf1), .Y(_3802_) );
	NAND2X1 NAND2X1_61 ( .A(_3802_), .B(_3801_), .Y(_3050__3_) );
	AND2X2 AND2X2_9 ( .A(_3795_), .B(_3718_), .Y(_3803_) );
	INVX1 INVX1_21 ( .A(micro_hash_synth_2_x_4_), .Y(_3804_) );
	NOR2X1 NOR2X1_19 ( .A(_3434_), .B(_3804_), .Y(_3805_) );
	NOR2X1 NOR2X1_20 ( .A(micro_hash_synth_2_k_4_), .B(micro_hash_synth_2_x_4_), .Y(_3806_) );
	NOR2X1 NOR2X1_21 ( .A(_3806_), .B(_3805_), .Y(_3807_) );
	NOR2X1 NOR2X1_22 ( .A(micro_hash_synth_2_W_29__4_), .B(_4733__bF_buf1), .Y(_3808_) );
	OAI21X1 OAI21X1_38 ( .A(concatenador_counter_2d_0_bF_buf6), .B(micro_hash_synth_2_W_28__4_), .C(concatenador_counter_2d_1_bF_buf4), .Y(_3809_) );
	NOR2X1 NOR2X1_23 ( .A(concatenador_counter_2d_0_bF_buf5), .B(micro_hash_synth_2_W_30__4_), .Y(_3810_) );
	OAI21X1 OAI21X1_39 ( .A(_4733__bF_buf0), .B(micro_hash_synth_2_W_31__4_), .C(_3439__bF_buf0), .Y(_3811_) );
	OAI22X1 OAI22X1_15 ( .A(_3808_), .B(_3809_), .C(_3811_), .D(_3810_), .Y(_3812_) );
	INVX1 INVX1_22 ( .A(micro_hash_synth_2_W_24__4_), .Y(_3813_) );
	NAND2X1 NAND2X1_62 ( .A(concatenador_counter_2d_0_bF_buf4), .B(micro_hash_synth_2_W_25__4_), .Y(_3814_) );
	OAI21X1 OAI21X1_40 ( .A(_3813_), .B(concatenador_counter_2d_0_bF_buf3), .C(_3814_), .Y(_3815_) );
	NAND2X1 NAND2X1_63 ( .A(_3440__bF_buf3), .B(_3815_), .Y(_3816_) );
	NAND2X1 NAND2X1_64 ( .A(concatenador_counter_2d_0_bF_buf2), .B(micro_hash_synth_2_W_27__4_), .Y(_3817_) );
	OAI21X1 OAI21X1_41 ( .A(_4756_), .B(concatenador_counter_2d_0_bF_buf1), .C(_3817_), .Y(_3818_) );
	NAND2X1 NAND2X1_65 ( .A(_3442__bF_buf1), .B(_3818_), .Y(_3819_) );
	NAND3X1 NAND3X1_32 ( .A(_3489__bF_buf3), .B(_3816_), .C(_3819_), .Y(_3820_) );
	AOI21X1 AOI21X1_24 ( .A(_3443__bF_buf1), .B(_3812_), .C(_3820_), .Y(_3821_) );
	NOR2X1 NOR2X1_24 ( .A(micro_hash_synth_2_W_13__4_), .B(_4733__bF_buf7), .Y(_3822_) );
	OAI21X1 OAI21X1_42 ( .A(concatenador_counter_2d_0_bF_buf0), .B(micro_hash_synth_2_W_12__4_), .C(concatenador_counter_2d_1_bF_buf3), .Y(_3823_) );
	NOR2X1 NOR2X1_25 ( .A(concatenador_counter_2d_0_bF_buf12), .B(micro_hash_synth_2_W_14__4_), .Y(_3824_) );
	OAI21X1 OAI21X1_43 ( .A(_4733__bF_buf6), .B(micro_hash_synth_2_W_15__4_), .C(_3439__bF_buf3), .Y(_3825_) );
	OAI22X1 OAI22X1_16 ( .A(_3822_), .B(_3823_), .C(_3825_), .D(_3824_), .Y(_3826_) );
	INVX1 INVX1_23 ( .A(micro_hash_synth_2_W_10__4_), .Y(_3827_) );
	NAND2X1 NAND2X1_66 ( .A(concatenador_counter_2d_0_bF_buf11), .B(micro_hash_synth_2_W_11__4_), .Y(_3828_) );
	OAI21X1 OAI21X1_44 ( .A(_3827_), .B(concatenador_counter_2d_0_bF_buf10), .C(_3828_), .Y(_3829_) );
	NAND2X1 NAND2X1_67 ( .A(_3442__bF_buf0), .B(_3829_), .Y(_3830_) );
	NAND2X1 NAND2X1_68 ( .A(concatenador_counter_2d_0_bF_buf9), .B(micro_hash_synth_2_W_9__4_), .Y(_3831_) );
	OAI21X1 OAI21X1_45 ( .A(_4808_), .B(concatenador_counter_2d_0_bF_buf8), .C(_3831_), .Y(_3832_) );
	NAND2X1 NAND2X1_69 ( .A(_3440__bF_buf2), .B(_3832_), .Y(_3833_) );
	NAND3X1 NAND3X1_33 ( .A(_3489__bF_buf2), .B(_3830_), .C(_3833_), .Y(_3834_) );
	AOI21X1 AOI21X1_25 ( .A(_3443__bF_buf0), .B(_3826_), .C(_3834_), .Y(_3835_) );
	NOR2X1 NOR2X1_26 ( .A(micro_hash_synth_2_W_21__4_), .B(_4733__bF_buf5), .Y(_3836_) );
	OAI21X1 OAI21X1_46 ( .A(concatenador_counter_2d_0_bF_buf7), .B(micro_hash_synth_2_W_20__4_), .C(concatenador_counter_2d_1_bF_buf2), .Y(_3837_) );
	MUX2X1 MUX2X1_5 ( .A(micro_hash_synth_2_W_23__4_), .B(micro_hash_synth_2_W_22__4_), .S(concatenador_counter_2d_0_bF_buf6), .Y(_3838_) );
	OAI22X1 OAI22X1_17 ( .A(_3838_), .B(concatenador_counter_2d_1_bF_buf1), .C(_3836_), .D(_3837_), .Y(_3839_) );
	AND2X2 AND2X2_10 ( .A(_3839_), .B(_3443__bF_buf5), .Y(_3840_) );
	INVX1 INVX1_24 ( .A(micro_hash_synth_2_W_18__4_), .Y(_3841_) );
	NAND2X1 NAND2X1_70 ( .A(concatenador_counter_2d_0_bF_buf5), .B(micro_hash_synth_2_W_19__4_), .Y(_3842_) );
	OAI21X1 OAI21X1_47 ( .A(_3841_), .B(concatenador_counter_2d_0_bF_buf4), .C(_3842_), .Y(_3843_) );
	NAND2X1 NAND2X1_71 ( .A(_3442__bF_buf4), .B(_3843_), .Y(_3844_) );
	INVX1 INVX1_25 ( .A(micro_hash_synth_2_W_16__4_), .Y(_3845_) );
	NAND2X1 NAND2X1_72 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_17__4_), .Y(_3846_) );
	OAI21X1 OAI21X1_48 ( .A(_3845_), .B(concatenador_counter_2d_0_bF_buf2), .C(_3846_), .Y(_3847_) );
	NAND2X1 NAND2X1_73 ( .A(_3440__bF_buf1), .B(_3847_), .Y(_3848_) );
	NAND3X1 NAND3X1_34 ( .A(_3453__bF_buf1), .B(_3844_), .C(_3848_), .Y(_3849_) );
	OAI21X1 OAI21X1_49 ( .A(_3840_), .B(_3849_), .C(_3460_), .Y(_3850_) );
	NOR2X1 NOR2X1_27 ( .A(micro_hash_synth_2_W_5__4_), .B(_4733__bF_buf4), .Y(_3851_) );
	OAI21X1 OAI21X1_50 ( .A(concatenador_counter_2d_0_bF_buf1), .B(micro_hash_synth_2_W_4__4_), .C(concatenador_counter_2d_1_bF_buf0), .Y(_3852_) );
	MUX2X1 MUX2X1_6 ( .A(micro_hash_synth_2_W_7__4_), .B(micro_hash_synth_2_W_6__4_), .S(concatenador_counter_2d_0_bF_buf0), .Y(_3853_) );
	OAI22X1 OAI22X1_18 ( .A(_3853_), .B(concatenador_counter_2d_1_bF_buf6), .C(_3851_), .D(_3852_), .Y(_3854_) );
	AND2X2 AND2X2_11 ( .A(_3854_), .B(_3443__bF_buf4), .Y(_3855_) );
	NAND2X1 NAND2X1_74 ( .A(concatenador_counter_2d_0_bF_buf12), .B(micro_hash_synth_2_W_1__4_), .Y(_3856_) );
	OAI21X1 OAI21X1_51 ( .A(_4845_), .B(concatenador_counter_2d_0_bF_buf11), .C(_3856_), .Y(_3857_) );
	NAND2X1 NAND2X1_75 ( .A(_3440__bF_buf0), .B(_3857_), .Y(_3858_) );
	NAND2X1 NAND2X1_76 ( .A(concatenador_counter_2d_0_bF_buf10), .B(micro_hash_synth_2_W_3__4_), .Y(_3859_) );
	OAI21X1 OAI21X1_52 ( .A(_4853_), .B(concatenador_counter_2d_0_bF_buf9), .C(_3859_), .Y(_3860_) );
	NAND2X1 NAND2X1_77 ( .A(_3442__bF_buf3), .B(_3860_), .Y(_3861_) );
	NAND3X1 NAND3X1_35 ( .A(_3453__bF_buf0), .B(_3858_), .C(_3861_), .Y(_3862_) );
	OAI21X1 OAI21X1_53 ( .A(_3855_), .B(_3862_), .C(_3490_), .Y(_3863_) );
	OAI22X1 OAI22X1_19 ( .A(_3850_), .B(_3821_), .C(_3835_), .D(_3863_), .Y(_3864_) );
	NOR2X1 NOR2X1_28 ( .A(_3807_), .B(_3864_), .Y(_3865_) );
	INVX1 INVX1_26 ( .A(_3807_), .Y(_3866_) );
	NAND2X1 NAND2X1_78 ( .A(_3443__bF_buf3), .B(_3812_), .Y(_3867_) );
	AND2X2 AND2X2_12 ( .A(_3816_), .B(_3819_), .Y(_3868_) );
	AOI21X1 AOI21X1_26 ( .A(_3867_), .B(_3868_), .C(_3453__bF_buf3), .Y(_3869_) );
	NAND2X1 NAND2X1_79 ( .A(_3443__bF_buf2), .B(_3839_), .Y(_3870_) );
	AND2X2 AND2X2_13 ( .A(_3844_), .B(_3848_), .Y(_3871_) );
	AOI21X1 AOI21X1_27 ( .A(_3870_), .B(_3871_), .C(_3489__bF_buf1), .Y(_3872_) );
	OAI21X1 OAI21X1_54 ( .A(_3869_), .B(_3872_), .C(_3460_), .Y(_3873_) );
	NAND2X1 NAND2X1_80 ( .A(_3443__bF_buf1), .B(_3826_), .Y(_3874_) );
	AND2X2 AND2X2_14 ( .A(_3830_), .B(_3833_), .Y(_3875_) );
	AOI21X1 AOI21X1_28 ( .A(_3874_), .B(_3875_), .C(_3453__bF_buf2), .Y(_3876_) );
	NAND2X1 NAND2X1_81 ( .A(_3443__bF_buf0), .B(_3854_), .Y(_3877_) );
	AND2X2 AND2X2_15 ( .A(_3858_), .B(_3861_), .Y(_3878_) );
	AOI21X1 AOI21X1_29 ( .A(_3877_), .B(_3878_), .C(_3489__bF_buf0), .Y(_3879_) );
	OAI21X1 OAI21X1_55 ( .A(_3876_), .B(_3879_), .C(_3490_), .Y(_3880_) );
	AOI21X1 AOI21X1_30 ( .A(_3873_), .B(_3880_), .C(_3866_), .Y(_3881_) );
	OAI21X1 OAI21X1_56 ( .A(_3865_), .B(_3881_), .C(_3803_), .Y(_3882_) );
	OAI21X1 OAI21X1_57 ( .A(_3429_), .B(_3719_), .C(_3795_), .Y(_3883_) );
	NOR2X1 NOR2X1_29 ( .A(_3881_), .B(_3865_), .Y(_3884_) );
	NAND2X1 NAND2X1_82 ( .A(_3883_), .B(_3884_), .Y(_3885_) );
	NAND2X1 NAND2X1_83 ( .A(_3885_), .B(_3882_), .Y(_3886_) );
	OAI22X1 OAI22X1_20 ( .A(_3704_), .B(_3714_), .C(_3796_), .D(_3717_), .Y(_3887_) );
	OAI21X1 OAI21X1_58 ( .A(_3710_), .B(_3887_), .C(_3797_), .Y(_3888_) );
	AND2X2 AND2X2_16 ( .A(_3888_), .B(_3886_), .Y(_3889_) );
	OAI21X1 OAI21X1_59 ( .A(_3888_), .B(_3886_), .C(_3603_), .Y(_3890_) );
	AOI21X1 AOI21X1_31 ( .A(micro_hash_synth_2_c_4_), .B(_3436_), .C(_3332__bF_buf0), .Y(_3891_) );
	OAI21X1 OAI21X1_60 ( .A(_3889_), .B(_3890_), .C(_3891_), .Y(_3050__4_) );
	OAI21X1 OAI21X1_61 ( .A(_3888_), .B(_3886_), .C(_3885_), .Y(_3892_) );
	XOR2X1 XOR2X1_1 ( .A(micro_hash_synth_2_k_5_), .B(micro_hash_synth_2_x_5_), .Y(_3893_) );
	MUX2X1 MUX2X1_7 ( .A(micro_hash_synth_2_W_21__5_), .B(micro_hash_synth_2_W_20__5_), .S(concatenador_counter_2d_0_bF_buf8), .Y(_3894_) );
	MUX2X1 MUX2X1_8 ( .A(micro_hash_synth_2_W_23__5_), .B(micro_hash_synth_2_W_22__5_), .S(concatenador_counter_2d_0_bF_buf7), .Y(_3895_) );
	MUX2X1 MUX2X1_9 ( .A(_3895_), .B(_3894_), .S(_3439__bF_buf2), .Y(_3896_) );
	AND2X2 AND2X2_17 ( .A(_3896_), .B(_3443__bF_buf5), .Y(_3897_) );
	INVX1 INVX1_27 ( .A(micro_hash_synth_2_W_18__5_), .Y(_3898_) );
	NAND2X1 NAND2X1_84 ( .A(concatenador_counter_2d_0_bF_buf6), .B(micro_hash_synth_2_W_19__5_), .Y(_3899_) );
	OAI21X1 OAI21X1_62 ( .A(_3898_), .B(concatenador_counter_2d_0_bF_buf5), .C(_3899_), .Y(_3900_) );
	NAND2X1 NAND2X1_85 ( .A(_3442__bF_buf2), .B(_3900_), .Y(_3901_) );
	INVX1 INVX1_28 ( .A(micro_hash_synth_2_W_16__5_), .Y(_3902_) );
	NAND2X1 NAND2X1_86 ( .A(concatenador_counter_2d_0_bF_buf4), .B(micro_hash_synth_2_W_17__5_), .Y(_3903_) );
	OAI21X1 OAI21X1_63 ( .A(_3902_), .B(concatenador_counter_2d_0_bF_buf3), .C(_3903_), .Y(_3904_) );
	NAND2X1 NAND2X1_87 ( .A(_3440__bF_buf4), .B(_3904_), .Y(_3905_) );
	NAND3X1 NAND3X1_36 ( .A(_3453__bF_buf1), .B(_3901_), .C(_3905_), .Y(_3906_) );
	NOR2X1 NOR2X1_30 ( .A(micro_hash_synth_2_W_29__5_), .B(_4733__bF_buf3), .Y(_3907_) );
	OAI21X1 OAI21X1_64 ( .A(concatenador_counter_2d_0_bF_buf2), .B(micro_hash_synth_2_W_28__5_), .C(concatenador_counter_2d_1_bF_buf5), .Y(_3908_) );
	MUX2X1 MUX2X1_10 ( .A(micro_hash_synth_2_W_31__5_), .B(micro_hash_synth_2_W_30__5_), .S(concatenador_counter_2d_0_bF_buf1), .Y(_3909_) );
	OAI22X1 OAI22X1_21 ( .A(_3909_), .B(concatenador_counter_2d_1_bF_buf4), .C(_3907_), .D(_3908_), .Y(_3910_) );
	AND2X2 AND2X2_18 ( .A(_3910_), .B(_3443__bF_buf4), .Y(_3911_) );
	NAND2X1 NAND2X1_88 ( .A(concatenador_counter_2d_0_bF_buf0), .B(micro_hash_synth_2_W_27__5_), .Y(_3912_) );
	OAI21X1 OAI21X1_65 ( .A(_4759_), .B(concatenador_counter_2d_0_bF_buf12), .C(_3912_), .Y(_3913_) );
	NAND2X1 NAND2X1_89 ( .A(_3442__bF_buf1), .B(_3913_), .Y(_3914_) );
	INVX1 INVX1_29 ( .A(micro_hash_synth_2_W_24__5_), .Y(_3915_) );
	NAND2X1 NAND2X1_90 ( .A(concatenador_counter_2d_0_bF_buf11), .B(micro_hash_synth_2_W_25__5_), .Y(_3916_) );
	OAI21X1 OAI21X1_66 ( .A(_3915_), .B(concatenador_counter_2d_0_bF_buf10), .C(_3916_), .Y(_3917_) );
	NAND2X1 NAND2X1_91 ( .A(_3440__bF_buf3), .B(_3917_), .Y(_3918_) );
	NAND3X1 NAND3X1_37 ( .A(_3489__bF_buf3), .B(_3914_), .C(_3918_), .Y(_3919_) );
	OAI22X1 OAI22X1_22 ( .A(_3897_), .B(_3906_), .C(_3911_), .D(_3919_), .Y(_3920_) );
	NAND2X1 NAND2X1_92 ( .A(_3460_), .B(_3920_), .Y(_3921_) );
	MUX2X1 MUX2X1_11 ( .A(micro_hash_synth_2_W_13__5_), .B(micro_hash_synth_2_W_12__5_), .S(concatenador_counter_2d_0_bF_buf9), .Y(_3922_) );
	MUX2X1 MUX2X1_12 ( .A(micro_hash_synth_2_W_15__5_), .B(micro_hash_synth_2_W_14__5_), .S(concatenador_counter_2d_0_bF_buf8), .Y(_3923_) );
	MUX2X1 MUX2X1_13 ( .A(_3923_), .B(_3922_), .S(_3439__bF_buf1), .Y(_3924_) );
	AND2X2 AND2X2_19 ( .A(_3924_), .B(_3443__bF_buf3), .Y(_3925_) );
	NAND2X1 NAND2X1_93 ( .A(concatenador_counter_2d_0_bF_buf7), .B(micro_hash_synth_2_W_9__5_), .Y(_3926_) );
	OAI21X1 OAI21X1_67 ( .A(_4810_), .B(concatenador_counter_2d_0_bF_buf6), .C(_3926_), .Y(_3927_) );
	NAND2X1 NAND2X1_94 ( .A(_3440__bF_buf2), .B(_3927_), .Y(_3928_) );
	INVX1 INVX1_30 ( .A(micro_hash_synth_2_W_10__5_), .Y(_3929_) );
	NAND2X1 NAND2X1_95 ( .A(concatenador_counter_2d_0_bF_buf5), .B(micro_hash_synth_2_W_11__5_), .Y(_3930_) );
	OAI21X1 OAI21X1_68 ( .A(_3929_), .B(concatenador_counter_2d_0_bF_buf4), .C(_3930_), .Y(_3931_) );
	NAND2X1 NAND2X1_96 ( .A(_3442__bF_buf0), .B(_3931_), .Y(_3932_) );
	NAND3X1 NAND3X1_38 ( .A(_3489__bF_buf2), .B(_3928_), .C(_3932_), .Y(_3933_) );
	NOR2X1 NOR2X1_31 ( .A(micro_hash_synth_2_W_5__5_), .B(_4733__bF_buf2), .Y(_3934_) );
	OAI21X1 OAI21X1_69 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_4__5_), .C(concatenador_counter_2d_1_bF_buf3), .Y(_3935_) );
	MUX2X1 MUX2X1_14 ( .A(micro_hash_synth_2_W_7__5_), .B(micro_hash_synth_2_W_6__5_), .S(concatenador_counter_2d_0_bF_buf2), .Y(_3936_) );
	OAI22X1 OAI22X1_23 ( .A(_3936_), .B(concatenador_counter_2d_1_bF_buf2), .C(_3934_), .D(_3935_), .Y(_3937_) );
	AND2X2 AND2X2_20 ( .A(_3937_), .B(_3443__bF_buf2), .Y(_3938_) );
	NAND2X1 NAND2X1_97 ( .A(concatenador_counter_2d_0_bF_buf1), .B(micro_hash_synth_2_W_3__5_), .Y(_3939_) );
	OAI21X1 OAI21X1_70 ( .A(_4854_), .B(concatenador_counter_2d_0_bF_buf0), .C(_3939_), .Y(_3940_) );
	NAND2X1 NAND2X1_98 ( .A(_3442__bF_buf4), .B(_3940_), .Y(_3941_) );
	NAND2X1 NAND2X1_99 ( .A(concatenador_counter_2d_0_bF_buf12), .B(micro_hash_synth_2_W_1__5_), .Y(_3942_) );
	OAI21X1 OAI21X1_71 ( .A(_4846_), .B(concatenador_counter_2d_0_bF_buf11), .C(_3942_), .Y(_3943_) );
	NAND2X1 NAND2X1_100 ( .A(_3440__bF_buf1), .B(_3943_), .Y(_3944_) );
	NAND3X1 NAND3X1_39 ( .A(_3453__bF_buf0), .B(_3941_), .C(_3944_), .Y(_3945_) );
	OAI22X1 OAI22X1_24 ( .A(_3925_), .B(_3933_), .C(_3938_), .D(_3945_), .Y(_3946_) );
	NAND2X1 NAND2X1_101 ( .A(_3490_), .B(_3946_), .Y(_3947_) );
	AOI21X1 AOI21X1_32 ( .A(_3921_), .B(_3947_), .C(_3893_), .Y(_3948_) );
	INVX1 INVX1_31 ( .A(_3893_), .Y(_3949_) );
	OR2X2 OR2X2_7 ( .A(_3897_), .B(_3906_), .Y(_3950_) );
	OR2X2 OR2X2_8 ( .A(_3911_), .B(_3919_), .Y(_3951_) );
	NAND3X1 NAND3X1_40 ( .A(_3460_), .B(_3950_), .C(_3951_), .Y(_3952_) );
	OR2X2 OR2X2_9 ( .A(_3925_), .B(_3933_), .Y(_3953_) );
	OR2X2 OR2X2_10 ( .A(_3938_), .B(_3945_), .Y(_3954_) );
	NAND3X1 NAND3X1_41 ( .A(_3490_), .B(_3953_), .C(_3954_), .Y(_3955_) );
	AOI21X1 AOI21X1_33 ( .A(_3952_), .B(_3955_), .C(_3949_), .Y(_3956_) );
	OAI22X1 OAI22X1_25 ( .A(_3805_), .B(_3881_), .C(_3956_), .D(_3948_), .Y(_3957_) );
	AOI21X1 AOI21X1_34 ( .A(_3807_), .B(_3864_), .C(_3805_), .Y(_3958_) );
	NAND3X1 NAND3X1_42 ( .A(_3949_), .B(_3952_), .C(_3955_), .Y(_3959_) );
	NAND3X1 NAND3X1_43 ( .A(_3893_), .B(_3921_), .C(_3947_), .Y(_3960_) );
	NAND3X1 NAND3X1_44 ( .A(_3959_), .B(_3960_), .C(_3958_), .Y(_3961_) );
	NAND2X1 NAND2X1_102 ( .A(_3961_), .B(_3957_), .Y(_3962_) );
	XNOR2X1 XNOR2X1_1 ( .A(_3892_), .B(_3962_), .Y(_3963_) );
	AOI21X1 AOI21X1_35 ( .A(micro_hash_synth_2_c_5_), .B(_3436_), .C(_3332__bF_buf3), .Y(_3964_) );
	OAI21X1 OAI21X1_72 ( .A(_3963_), .B(_3505_), .C(_3964_), .Y(_3050__5_) );
	NAND3X1 NAND3X1_45 ( .A(_3882_), .B(_3885_), .C(_3962_), .Y(_3965_) );
	AND2X2 AND2X2_21 ( .A(_3884_), .B(_3883_), .Y(_3966_) );
	NAND2X1 NAND2X1_103 ( .A(_3960_), .B(_3959_), .Y(_3967_) );
	NOR2X1 NOR2X1_32 ( .A(_3958_), .B(_3967_), .Y(_3968_) );
	AOI21X1 AOI21X1_36 ( .A(_3962_), .B(_3966_), .C(_3968_), .Y(_3969_) );
	OAI21X1 OAI21X1_73 ( .A(_3888_), .B(_3965_), .C(_3969_), .Y(_3970_) );
	AOI21X1 AOI21X1_37 ( .A(micro_hash_synth_2_k_5_), .B(micro_hash_synth_2_x_5_), .C(_3956_), .Y(_3971_) );
	INVX1 INVX1_32 ( .A(_3971_), .Y(_3972_) );
	AND2X2 AND2X2_22 ( .A(micro_hash_synth_2_k_6_), .B(micro_hash_synth_2_x_6_), .Y(_3973_) );
	NOR2X1 NOR2X1_33 ( .A(micro_hash_synth_2_k_6_), .B(micro_hash_synth_2_x_6_), .Y(_3974_) );
	NOR2X1 NOR2X1_34 ( .A(_3974_), .B(_3973_), .Y(_3975_) );
	INVX1 INVX1_33 ( .A(_3975_), .Y(_3976_) );
	NOR2X1 NOR2X1_35 ( .A(micro_hash_synth_2_W_21__6_), .B(_4733__bF_buf1), .Y(_3977_) );
	OAI21X1 OAI21X1_74 ( .A(concatenador_counter_2d_0_bF_buf10), .B(micro_hash_synth_2_W_20__6_), .C(concatenador_counter_2d_1_bF_buf1), .Y(_3978_) );
	AOI21X1 AOI21X1_38 ( .A(concatenador_counter_2d_0_bF_buf9), .B(_4764_), .C(concatenador_counter_2d_1_bF_buf0), .Y(_3979_) );
	OAI21X1 OAI21X1_75 ( .A(concatenador_counter_2d_0_bF_buf8), .B(micro_hash_synth_2_W_22__6_), .C(_3979_), .Y(_3980_) );
	OAI21X1 OAI21X1_76 ( .A(_3977_), .B(_3978_), .C(_3980_), .Y(_3981_) );
	INVX1 INVX1_34 ( .A(micro_hash_synth_2_W_18__6_), .Y(_3982_) );
	AOI21X1 AOI21X1_39 ( .A(_4733__bF_buf0), .B(_3982_), .C(_3468_), .Y(_3983_) );
	OAI21X1 OAI21X1_77 ( .A(_4733__bF_buf7), .B(micro_hash_synth_2_W_19__6_), .C(_3983_), .Y(_3984_) );
	INVX1 INVX1_35 ( .A(micro_hash_synth_2_W_16__6_), .Y(_3985_) );
	AOI21X1 AOI21X1_40 ( .A(_4733__bF_buf6), .B(_3985_), .C(_3467_), .Y(_3986_) );
	OAI21X1 OAI21X1_78 ( .A(_4733__bF_buf5), .B(micro_hash_synth_2_W_17__6_), .C(_3986_), .Y(_3987_) );
	NAND2X1 NAND2X1_104 ( .A(_3984_), .B(_3987_), .Y(_3988_) );
	AOI21X1 AOI21X1_41 ( .A(_3443__bF_buf1), .B(_3981_), .C(_3988_), .Y(_3989_) );
	NOR2X1 NOR2X1_36 ( .A(micro_hash_synth_2_W_29__6_), .B(_4733__bF_buf4), .Y(_3990_) );
	OAI21X1 OAI21X1_79 ( .A(concatenador_counter_2d_0_bF_buf7), .B(micro_hash_synth_2_W_28__6_), .C(concatenador_counter_2d_1_bF_buf6), .Y(_3991_) );
	NOR2X1 NOR2X1_37 ( .A(concatenador_counter_2d_0_bF_buf6), .B(micro_hash_synth_2_W_30__6_), .Y(_3992_) );
	OAI21X1 OAI21X1_80 ( .A(_4733__bF_buf3), .B(micro_hash_synth_2_W_31__6_), .C(_3439__bF_buf0), .Y(_3993_) );
	OAI22X1 OAI22X1_26 ( .A(_3990_), .B(_3991_), .C(_3993_), .D(_3992_), .Y(_3994_) );
	AND2X2 AND2X2_23 ( .A(_3994_), .B(_3443__bF_buf0), .Y(_3995_) );
	INVX1 INVX1_36 ( .A(micro_hash_synth_2_W_24__6_), .Y(_3996_) );
	AOI21X1 AOI21X1_42 ( .A(_4733__bF_buf2), .B(_3996_), .C(_3467_), .Y(_3997_) );
	OAI21X1 OAI21X1_81 ( .A(_4733__bF_buf1), .B(micro_hash_synth_2_W_25__6_), .C(_3997_), .Y(_3998_) );
	AOI21X1 AOI21X1_43 ( .A(_4733__bF_buf0), .B(_4762_), .C(_3468_), .Y(_3999_) );
	OAI21X1 OAI21X1_82 ( .A(_4733__bF_buf7), .B(micro_hash_synth_2_W_27__6_), .C(_3999_), .Y(_4000_) );
	NAND2X1 NAND2X1_105 ( .A(_3998_), .B(_4000_), .Y(_4001_) );
	OAI21X1 OAI21X1_83 ( .A(_4001_), .B(_3995_), .C(_3489__bF_buf1), .Y(_4002_) );
	OAI21X1 OAI21X1_84 ( .A(_3489__bF_buf0), .B(_3989_), .C(_4002_), .Y(_4003_) );
	NAND2X1 NAND2X1_106 ( .A(_3460_), .B(_4003_), .Y(_4004_) );
	NOR2X1 NOR2X1_38 ( .A(micro_hash_synth_2_W_13__6_), .B(_4733__bF_buf6), .Y(_4005_) );
	OAI21X1 OAI21X1_85 ( .A(concatenador_counter_2d_0_bF_buf5), .B(micro_hash_synth_2_W_12__6_), .C(concatenador_counter_2d_1_bF_buf5), .Y(_4006_) );
	INVX1 INVX1_37 ( .A(micro_hash_synth_2_W_15__6_), .Y(_4007_) );
	AOI21X1 AOI21X1_44 ( .A(concatenador_counter_2d_0_bF_buf4), .B(_4007_), .C(concatenador_counter_2d_1_bF_buf4), .Y(_4008_) );
	OAI21X1 OAI21X1_86 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_14__6_), .C(_4008_), .Y(_4009_) );
	OAI21X1 OAI21X1_87 ( .A(_4005_), .B(_4006_), .C(_4009_), .Y(_4010_) );
	AND2X2 AND2X2_24 ( .A(_4010_), .B(_3443__bF_buf5), .Y(_4011_) );
	INVX1 INVX1_38 ( .A(micro_hash_synth_2_W_9__6_), .Y(_4012_) );
	AOI21X1 AOI21X1_45 ( .A(concatenador_counter_2d_0_bF_buf2), .B(_4012_), .C(_3467_), .Y(_4013_) );
	OAI21X1 OAI21X1_88 ( .A(concatenador_counter_2d_0_bF_buf1), .B(micro_hash_synth_2_W_8__6_), .C(_4013_), .Y(_4014_) );
	INVX1 INVX1_39 ( .A(micro_hash_synth_2_W_10__6_), .Y(_4015_) );
	AOI21X1 AOI21X1_46 ( .A(_4733__bF_buf5), .B(_4015_), .C(_3468_), .Y(_4016_) );
	OAI21X1 OAI21X1_89 ( .A(_4733__bF_buf4), .B(micro_hash_synth_2_W_11__6_), .C(_4016_), .Y(_4017_) );
	NAND2X1 NAND2X1_107 ( .A(_4014_), .B(_4017_), .Y(_4018_) );
	OAI21X1 OAI21X1_90 ( .A(_4011_), .B(_4018_), .C(_3489__bF_buf3), .Y(_4019_) );
	NOR2X1 NOR2X1_39 ( .A(micro_hash_synth_2_W_5__6_), .B(_4733__bF_buf3), .Y(_4020_) );
	OAI21X1 OAI21X1_91 ( .A(concatenador_counter_2d_0_bF_buf0), .B(micro_hash_synth_2_W_4__6_), .C(concatenador_counter_2d_1_bF_buf3), .Y(_4021_) );
	INVX1 INVX1_40 ( .A(micro_hash_synth_2_W_7__6_), .Y(_4022_) );
	AOI21X1 AOI21X1_47 ( .A(concatenador_counter_2d_0_bF_buf12), .B(_4022_), .C(concatenador_counter_2d_1_bF_buf2), .Y(_4023_) );
	OAI21X1 OAI21X1_92 ( .A(concatenador_counter_2d_0_bF_buf11), .B(micro_hash_synth_2_W_6__6_), .C(_4023_), .Y(_4024_) );
	OAI21X1 OAI21X1_93 ( .A(_4020_), .B(_4021_), .C(_4024_), .Y(_4025_) );
	AND2X2 AND2X2_25 ( .A(_4025_), .B(_3443__bF_buf4), .Y(_4026_) );
	AOI21X1 AOI21X1_48 ( .A(concatenador_counter_2d_0_bF_buf10), .B(_4839_), .C(_3467_), .Y(_4027_) );
	OAI21X1 OAI21X1_94 ( .A(concatenador_counter_2d_0_bF_buf9), .B(micro_hash_synth_2_W_0__6_), .C(_4027_), .Y(_4028_) );
	AOI21X1 AOI21X1_49 ( .A(_4733__bF_buf2), .B(_4855_), .C(_3468_), .Y(_4029_) );
	OAI21X1 OAI21X1_95 ( .A(_4733__bF_buf1), .B(micro_hash_synth_2_W_3__6_), .C(_4029_), .Y(_4030_) );
	NAND2X1 NAND2X1_108 ( .A(_4028_), .B(_4030_), .Y(_4031_) );
	OAI21X1 OAI21X1_96 ( .A(_4026_), .B(_4031_), .C(_3453__bF_buf3), .Y(_4032_) );
	NAND2X1 NAND2X1_109 ( .A(_4019_), .B(_4032_), .Y(_4033_) );
	NAND2X1 NAND2X1_110 ( .A(_3490_), .B(_4033_), .Y(_4034_) );
	NAND3X1 NAND3X1_46 ( .A(_3976_), .B(_4004_), .C(_4034_), .Y(_4035_) );
	INVX1 INVX1_41 ( .A(_4035_), .Y(_4036_) );
	AOI21X1 AOI21X1_50 ( .A(_4004_), .B(_4034_), .C(_3976_), .Y(_4037_) );
	OAI21X1 OAI21X1_97 ( .A(_4036_), .B(_4037_), .C(_3972_), .Y(_4038_) );
	INVX1 INVX1_42 ( .A(_4037_), .Y(_4039_) );
	NAND3X1 NAND3X1_47 ( .A(_3971_), .B(_4035_), .C(_4039_), .Y(_4040_) );
	NAND2X1 NAND2X1_111 ( .A(_4038_), .B(_4040_), .Y(_4041_) );
	XNOR2X1 XNOR2X1_2 ( .A(_3970_), .B(_4041_), .Y(_4042_) );
	AOI21X1 AOI21X1_51 ( .A(micro_hash_synth_2_c_6_), .B(_3436_), .C(_3332__bF_buf2), .Y(_4043_) );
	OAI21X1 OAI21X1_98 ( .A(_4042_), .B(_3505_), .C(_4043_), .Y(_3050__6_) );
	NAND2X1 NAND2X1_112 ( .A(_4035_), .B(_4039_), .Y(_4044_) );
	NOR2X1 NOR2X1_40 ( .A(_3971_), .B(_4044_), .Y(_4045_) );
	AOI21X1 AOI21X1_52 ( .A(_4041_), .B(_3970_), .C(_4045_), .Y(_4046_) );
	NOR2X1 NOR2X1_41 ( .A(micro_hash_synth_2_W_21__7_), .B(_4733__bF_buf0), .Y(_4047_) );
	OAI21X1 OAI21X1_99 ( .A(concatenador_counter_2d_0_bF_buf8), .B(micro_hash_synth_2_W_20__7_), .C(concatenador_counter_2d_1_bF_buf1), .Y(_4048_) );
	AOI21X1 AOI21X1_53 ( .A(concatenador_counter_2d_0_bF_buf7), .B(_4769_), .C(concatenador_counter_2d_1_bF_buf0), .Y(_4049_) );
	OAI21X1 OAI21X1_100 ( .A(concatenador_counter_2d_0_bF_buf6), .B(micro_hash_synth_2_W_22__7_), .C(_4049_), .Y(_4050_) );
	OAI21X1 OAI21X1_101 ( .A(_4047_), .B(_4048_), .C(_4050_), .Y(_4051_) );
	INVX1 INVX1_43 ( .A(micro_hash_synth_2_W_18__7_), .Y(_4052_) );
	AOI21X1 AOI21X1_54 ( .A(_4733__bF_buf7), .B(_4052_), .C(_3468_), .Y(_4053_) );
	OAI21X1 OAI21X1_102 ( .A(_4733__bF_buf6), .B(micro_hash_synth_2_W_19__7_), .C(_4053_), .Y(_4054_) );
	NOR2X1 NOR2X1_42 ( .A(micro_hash_synth_2_W_17__7_), .B(_4733__bF_buf5), .Y(_4055_) );
	OAI21X1 OAI21X1_103 ( .A(concatenador_counter_2d_0_bF_buf5), .B(micro_hash_synth_2_W_16__7_), .C(_3440__bF_buf0), .Y(_4056_) );
	OAI21X1 OAI21X1_104 ( .A(_4055_), .B(_4056_), .C(_4054_), .Y(_4057_) );
	AOI21X1 AOI21X1_55 ( .A(_3443__bF_buf3), .B(_4051_), .C(_4057_), .Y(_4058_) );
	NAND2X1 NAND2X1_113 ( .A(_3453__bF_buf2), .B(_4058_), .Y(_4059_) );
	NOR2X1 NOR2X1_43 ( .A(micro_hash_synth_2_W_29__7_), .B(_4733__bF_buf4), .Y(_4060_) );
	OAI21X1 OAI21X1_105 ( .A(concatenador_counter_2d_0_bF_buf4), .B(micro_hash_synth_2_W_28__7_), .C(concatenador_counter_2d_1_bF_buf6), .Y(_4061_) );
	NOR2X1 NOR2X1_44 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_30__7_), .Y(_4062_) );
	OAI21X1 OAI21X1_106 ( .A(_4733__bF_buf3), .B(micro_hash_synth_2_W_31__7_), .C(_3439__bF_buf3), .Y(_4063_) );
	OAI22X1 OAI22X1_27 ( .A(_4060_), .B(_4061_), .C(_4063_), .D(_4062_), .Y(_4064_) );
	NAND2X1 NAND2X1_114 ( .A(_3443__bF_buf2), .B(_4064_), .Y(_4065_) );
	AOI21X1 AOI21X1_56 ( .A(_4733__bF_buf2), .B(_4767_), .C(_3468_), .Y(_4066_) );
	OAI21X1 OAI21X1_107 ( .A(_4733__bF_buf1), .B(micro_hash_synth_2_W_27__7_), .C(_4066_), .Y(_4067_) );
	INVX1 INVX1_44 ( .A(micro_hash_synth_2_W_24__7_), .Y(_4068_) );
	AOI21X1 AOI21X1_57 ( .A(_4733__bF_buf0), .B(_4068_), .C(_3467_), .Y(_4069_) );
	OAI21X1 OAI21X1_108 ( .A(_4733__bF_buf7), .B(micro_hash_synth_2_W_25__7_), .C(_4069_), .Y(_4070_) );
	NAND3X1 NAND3X1_48 ( .A(_4067_), .B(_4070_), .C(_4065_), .Y(_4071_) );
	OAI21X1 OAI21X1_109 ( .A(_3453__bF_buf1), .B(_4071_), .C(_4059_), .Y(_4072_) );
	NAND2X1 NAND2X1_115 ( .A(_3460_), .B(_4072_), .Y(_4073_) );
	NOR2X1 NOR2X1_45 ( .A(micro_hash_synth_2_W_13__7_), .B(_4733__bF_buf6), .Y(_4074_) );
	OAI21X1 OAI21X1_110 ( .A(concatenador_counter_2d_0_bF_buf2), .B(micro_hash_synth_2_W_12__7_), .C(concatenador_counter_2d_1_bF_buf5), .Y(_4075_) );
	INVX1 INVX1_45 ( .A(micro_hash_synth_2_W_15__7_), .Y(_4076_) );
	AOI21X1 AOI21X1_58 ( .A(concatenador_counter_2d_0_bF_buf1), .B(_4076_), .C(concatenador_counter_2d_1_bF_buf4), .Y(_4077_) );
	OAI21X1 OAI21X1_111 ( .A(concatenador_counter_2d_0_bF_buf0), .B(micro_hash_synth_2_W_14__7_), .C(_4077_), .Y(_4078_) );
	OAI21X1 OAI21X1_112 ( .A(_4074_), .B(_4075_), .C(_4078_), .Y(_4079_) );
	AOI21X1 AOI21X1_59 ( .A(_4733__bF_buf5), .B(_4814_), .C(_3467_), .Y(_4080_) );
	OAI21X1 OAI21X1_113 ( .A(_4733__bF_buf4), .B(micro_hash_synth_2_W_9__7_), .C(_4080_), .Y(_4081_) );
	NOR2X1 NOR2X1_46 ( .A(micro_hash_synth_2_W_11__7_), .B(_4733__bF_buf3), .Y(_4082_) );
	OAI21X1 OAI21X1_114 ( .A(concatenador_counter_2d_0_bF_buf12), .B(micro_hash_synth_2_W_10__7_), .C(_3442__bF_buf3), .Y(_4083_) );
	OAI21X1 OAI21X1_115 ( .A(_4082_), .B(_4083_), .C(_4081_), .Y(_4084_) );
	AOI21X1 AOI21X1_60 ( .A(_3443__bF_buf1), .B(_4079_), .C(_4084_), .Y(_4085_) );
	NAND2X1 NAND2X1_116 ( .A(_3489__bF_buf2), .B(_4085_), .Y(_4086_) );
	NOR2X1 NOR2X1_47 ( .A(micro_hash_synth_2_W_5__7_), .B(_4733__bF_buf2), .Y(_4087_) );
	OAI21X1 OAI21X1_116 ( .A(concatenador_counter_2d_0_bF_buf11), .B(micro_hash_synth_2_W_4__7_), .C(concatenador_counter_2d_1_bF_buf3), .Y(_4088_) );
	NOR2X1 NOR2X1_48 ( .A(_4088_), .B(_4087_), .Y(_4089_) );
	INVX1 INVX1_46 ( .A(micro_hash_synth_2_W_6__7_), .Y(_4090_) );
	OAI21X1 OAI21X1_117 ( .A(_4733__bF_buf1), .B(micro_hash_synth_2_W_7__7_), .C(_3439__bF_buf2), .Y(_4091_) );
	AOI21X1 AOI21X1_61 ( .A(_4733__bF_buf0), .B(_4090_), .C(_4091_), .Y(_4092_) );
	OAI21X1 OAI21X1_118 ( .A(_4092_), .B(_4089_), .C(_3443__bF_buf0), .Y(_4093_) );
	AOI21X1 AOI21X1_62 ( .A(_4733__bF_buf7), .B(_4848_), .C(_3467_), .Y(_4094_) );
	OAI21X1 OAI21X1_119 ( .A(_4733__bF_buf6), .B(micro_hash_synth_2_W_1__7_), .C(_4094_), .Y(_4095_) );
	AOI21X1 AOI21X1_63 ( .A(_4733__bF_buf5), .B(_4856_), .C(_3468_), .Y(_4096_) );
	OAI21X1 OAI21X1_120 ( .A(_4733__bF_buf4), .B(micro_hash_synth_2_W_3__7_), .C(_4096_), .Y(_4097_) );
	NAND3X1 NAND3X1_49 ( .A(_4095_), .B(_4097_), .C(_4093_), .Y(_4098_) );
	OAI21X1 OAI21X1_121 ( .A(_3489__bF_buf1), .B(_4098_), .C(_4086_), .Y(_4099_) );
	NAND2X1 NAND2X1_117 ( .A(_3490_), .B(_4099_), .Y(_4100_) );
	AND2X2 AND2X2_26 ( .A(_4073_), .B(_4100_), .Y(_4101_) );
	XOR2X1 XOR2X1_2 ( .A(micro_hash_synth_2_k_7_), .B(micro_hash_synth_2_x_7_), .Y(_4102_) );
	INVX1 INVX1_47 ( .A(_4102_), .Y(_4103_) );
	NOR2X1 NOR2X1_49 ( .A(_4103_), .B(_4101_), .Y(_4104_) );
	NAND2X1 NAND2X1_118 ( .A(_4073_), .B(_4100_), .Y(_4105_) );
	NOR2X1 NOR2X1_50 ( .A(_4102_), .B(_4105_), .Y(_4106_) );
	OAI22X1 OAI22X1_28 ( .A(_3973_), .B(_4037_), .C(_4104_), .D(_4106_), .Y(_4107_) );
	NOR2X1 NOR2X1_51 ( .A(_3973_), .B(_4037_), .Y(_4108_) );
	NOR2X1 NOR2X1_52 ( .A(_4102_), .B(_4101_), .Y(_4109_) );
	NOR2X1 NOR2X1_53 ( .A(_4103_), .B(_4105_), .Y(_4110_) );
	OAI21X1 OAI21X1_122 ( .A(_4109_), .B(_4110_), .C(_4108_), .Y(_4111_) );
	NAND2X1 NAND2X1_119 ( .A(_4111_), .B(_4107_), .Y(_4112_) );
	XNOR2X1 XNOR2X1_3 ( .A(_4046_), .B(_4112_), .Y(_4113_) );
	AOI21X1 AOI21X1_64 ( .A(micro_hash_synth_2_c_7_), .B(_3436_), .C(_3332__bF_buf1), .Y(_4114_) );
	OAI21X1 OAI21X1_123 ( .A(_4113_), .B(_3505_), .C(_4114_), .Y(_3050__7_) );
	OAI21X1 OAI21X1_124 ( .A(_3322_), .B(_3424__bF_buf3), .C(_3333__bF_buf3), .Y(_3049__0_) );
	NOR2X1 NOR2X1_54 ( .A(_3325_), .B(_3426_), .Y(_3049__1_) );
	INVX1 INVX1_48 ( .A(micro_hash_synth_2_b_2_), .Y(_4115_) );
	NOR2X1 NOR2X1_55 ( .A(_4115_), .B(_3426_), .Y(_3049__2_) );
	OAI21X1 OAI21X1_125 ( .A(_3343_), .B(_3424__bF_buf2), .C(_3333__bF_buf2), .Y(_3049__3_) );
	OAI21X1 OAI21X1_126 ( .A(micro_hash_synth_2_b_4_), .B(_3424__bF_buf1), .C(_3333__bF_buf1), .Y(_4116_) );
	AOI21X1 AOI21X1_65 ( .A(_3438_), .B(_3603_), .C(_4116_), .Y(_3049__4_) );
	INVX1 INVX1_49 ( .A(micro_hash_synth_2_c_1_), .Y(_4117_) );
	OAI21X1 OAI21X1_127 ( .A(micro_hash_synth_2_b_5_), .B(_3424__bF_buf0), .C(_3333__bF_buf0), .Y(_4118_) );
	AOI21X1 AOI21X1_66 ( .A(_4117_), .B(_3603_), .C(_4118_), .Y(_3049__5_) );
	INVX1 INVX1_50 ( .A(micro_hash_synth_2_c_2_), .Y(_4119_) );
	OAI21X1 OAI21X1_128 ( .A(micro_hash_synth_2_b_6_), .B(_3424__bF_buf3), .C(_3333__bF_buf3), .Y(_4120_) );
	AOI21X1 AOI21X1_67 ( .A(_4119_), .B(_3603_), .C(_4120_), .Y(_3049__6_) );
	INVX1 INVX1_51 ( .A(micro_hash_synth_2_b_7_), .Y(_4121_) );
	NOR2X1 NOR2X1_56 ( .A(micro_hash_synth_2_c_3_), .B(_3436_), .Y(_4122_) );
	AOI22X1 AOI22X1_1 ( .A(_4121_), .B(_3425_), .C(_4122_), .D(_3333__bF_buf2), .Y(_3049__7_) );
	XNOR2X1 XNOR2X1_4 ( .A(micro_hash_synth_2_b_0_), .B(micro_hash_synth_2_c_0_), .Y(_4123_) );
	AOI21X1 AOI21X1_68 ( .A(micro_hash_synth_2_a_0_), .B(_3436_), .C(_3332__bF_buf0), .Y(_4124_) );
	OAI21X1 OAI21X1_129 ( .A(_3505_), .B(_4123_), .C(_4124_), .Y(_3048__0_) );
	NOR2X1 NOR2X1_57 ( .A(micro_hash_synth_2_b_1_), .B(_4117_), .Y(_4125_) );
	NOR2X1 NOR2X1_58 ( .A(micro_hash_synth_2_c_1_), .B(_3325_), .Y(_4126_) );
	OAI21X1 OAI21X1_130 ( .A(_4125_), .B(_4126_), .C(_3603_), .Y(_4127_) );
	OAI22X1 OAI22X1_29 ( .A(_3378_), .B(_3426_), .C(_4127_), .D(_4832__bF_buf5), .Y(_3048__1_) );
	INVX1 INVX1_52 ( .A(micro_hash_synth_2_a_2_), .Y(_4128_) );
	NOR2X1 NOR2X1_59 ( .A(micro_hash_synth_2_b_2_), .B(_4119_), .Y(_4129_) );
	NOR2X1 NOR2X1_60 ( .A(micro_hash_synth_2_c_2_), .B(_4115_), .Y(_4130_) );
	OAI21X1 OAI21X1_131 ( .A(_4129_), .B(_4130_), .C(_3603_), .Y(_4131_) );
	OAI22X1 OAI22X1_30 ( .A(_4128_), .B(_3426_), .C(_4131_), .D(_4832__bF_buf4), .Y(_3048__2_) );
	NAND2X1 NAND2X1_120 ( .A(micro_hash_synth_2_a_3_), .B(_3425_), .Y(_4132_) );
	INVX1 INVX1_53 ( .A(micro_hash_synth_2_c_3_), .Y(_4133_) );
	NOR2X1 NOR2X1_61 ( .A(micro_hash_synth_2_b_3_), .B(_4133_), .Y(_4134_) );
	NOR2X1 NOR2X1_62 ( .A(micro_hash_synth_2_c_3_), .B(_3343_), .Y(_4135_) );
	OAI21X1 OAI21X1_132 ( .A(_4134_), .B(_4135_), .C(_3603_), .Y(_4136_) );
	OAI21X1 OAI21X1_133 ( .A(_4136_), .B(_4832__bF_buf3), .C(_4132_), .Y(_3048__3_) );
	INVX1 INVX1_54 ( .A(micro_hash_synth_2_a_4_), .Y(_4137_) );
	INVX1 INVX1_55 ( .A(micro_hash_synth_2_c_4_), .Y(_4138_) );
	NOR2X1 NOR2X1_63 ( .A(micro_hash_synth_2_b_4_), .B(_4138_), .Y(_4139_) );
	INVX1 INVX1_56 ( .A(micro_hash_synth_2_b_4_), .Y(_4140_) );
	NOR2X1 NOR2X1_64 ( .A(micro_hash_synth_2_c_4_), .B(_4140_), .Y(_4141_) );
	OAI21X1 OAI21X1_134 ( .A(_4139_), .B(_4141_), .C(_3603_), .Y(_4142_) );
	OAI22X1 OAI22X1_31 ( .A(_4137_), .B(_3426_), .C(_4142_), .D(_4832__bF_buf2), .Y(_3048__4_) );
	NAND2X1 NAND2X1_121 ( .A(micro_hash_synth_2_a_5_), .B(_3425_), .Y(_4143_) );
	INVX1 INVX1_57 ( .A(micro_hash_synth_2_c_5_), .Y(_4144_) );
	NOR2X1 NOR2X1_65 ( .A(micro_hash_synth_2_b_5_), .B(_4144_), .Y(_4145_) );
	AND2X2 AND2X2_27 ( .A(_4144_), .B(micro_hash_synth_2_b_5_), .Y(_4146_) );
	OAI21X1 OAI21X1_135 ( .A(_4145_), .B(_4146_), .C(_3603_), .Y(_4147_) );
	OAI21X1 OAI21X1_136 ( .A(_4147_), .B(_4832__bF_buf1), .C(_4143_), .Y(_3048__5_) );
	INVX1 INVX1_58 ( .A(micro_hash_synth_2_c_6_), .Y(_4148_) );
	NOR2X1 NOR2X1_66 ( .A(micro_hash_synth_2_b_6_), .B(_4148_), .Y(_4149_) );
	AND2X2 AND2X2_28 ( .A(_4148_), .B(micro_hash_synth_2_b_6_), .Y(_4150_) );
	OAI21X1 OAI21X1_137 ( .A(_4149_), .B(_4150_), .C(_3603_), .Y(_4151_) );
	OAI22X1 OAI22X1_32 ( .A(_3418_), .B(_3426_), .C(_4151_), .D(_4832__bF_buf0), .Y(_3048__6_) );
	INVX1 INVX1_59 ( .A(micro_hash_synth_2_a_7_), .Y(_4152_) );
	AND2X2 AND2X2_29 ( .A(_4121_), .B(micro_hash_synth_2_c_7_), .Y(_4153_) );
	NOR2X1 NOR2X1_67 ( .A(micro_hash_synth_2_c_7_), .B(_4121_), .Y(_4154_) );
	OAI21X1 OAI21X1_138 ( .A(_4153_), .B(_4154_), .C(_3603_), .Y(_4155_) );
	OAI22X1 OAI22X1_33 ( .A(_4152_), .B(_3426_), .C(_4155_), .D(_4832__bF_buf5), .Y(_3048__7_) );
	XNOR2X1 XNOR2X1_5 ( .A(micro_hash_synth_2_c_0_), .B(Hhash_synth2_16_), .Y(_4156_) );
	NAND2X1 NAND2X1_122 ( .A(Hhash_synth2_16_), .B(_3333__bF_buf1), .Y(_4157_) );
	AOI22X1 AOI22X1_2 ( .A(_3316__bF_buf3), .B(_4156_), .C(_3320_), .D(_4157_), .Y(_3047__16_) );
	INVX1 INVX1_60 ( .A(Hhash_synth2_17_), .Y(_4158_) );
	NOR2X1 NOR2X1_68 ( .A(_4117_), .B(_4158_), .Y(_4159_) );
	NOR2X1 NOR2X1_69 ( .A(micro_hash_synth_2_c_1_), .B(Hhash_synth2_17_), .Y(_4160_) );
	NOR2X1 NOR2X1_70 ( .A(_4160_), .B(_4159_), .Y(_4161_) );
	NAND3X1 NAND3X1_50 ( .A(micro_hash_synth_2_c_0_), .B(Hhash_synth2_16_), .C(_4161_), .Y(_4162_) );
	NAND2X1 NAND2X1_123 ( .A(micro_hash_synth_2_c_0_), .B(Hhash_synth2_16_), .Y(_4163_) );
	OAI21X1 OAI21X1_139 ( .A(_4159_), .B(_4160_), .C(_4163_), .Y(_4164_) );
	NAND3X1 NAND3X1_51 ( .A(_4162_), .B(_4164_), .C(_3316__bF_buf2), .Y(_4165_) );
	OAI21X1 OAI21X1_140 ( .A(_4738_), .B(Hhash_synth2_17_), .C(_3317_), .Y(_4166_) );
	NAND3X1 NAND3X1_52 ( .A(reset_L_bF_buf49), .B(_4165_), .C(_4166_), .Y(_3047__17_) );
	OAI21X1 OAI21X1_141 ( .A(Hhash_synth2_18_), .B(_3332__bF_buf3), .C(_3320_), .Y(_4167_) );
	OAI21X1 OAI21X1_142 ( .A(_4117_), .B(_4158_), .C(_4162_), .Y(_4168_) );
	INVX1 INVX1_61 ( .A(Hhash_synth2_18_), .Y(_4169_) );
	NOR2X1 NOR2X1_71 ( .A(_4119_), .B(_4169_), .Y(_4170_) );
	NOR2X1 NOR2X1_72 ( .A(micro_hash_synth_2_c_2_), .B(Hhash_synth2_18_), .Y(_4171_) );
	NOR2X1 NOR2X1_73 ( .A(_4171_), .B(_4170_), .Y(_4172_) );
	NOR2X1 NOR2X1_74 ( .A(_4172_), .B(_4168_), .Y(_4173_) );
	NAND2X1 NAND2X1_124 ( .A(_4172_), .B(_4168_), .Y(_4174_) );
	NAND2X1 NAND2X1_125 ( .A(_4174_), .B(_3316__bF_buf1), .Y(_4175_) );
	OAI21X1 OAI21X1_143 ( .A(_4175_), .B(_4173_), .C(_4167_), .Y(_3047__18_) );
	AOI21X1 AOI21X1_69 ( .A(_4172_), .B(_4168_), .C(_4170_), .Y(_4176_) );
	INVX1 INVX1_62 ( .A(Hhash_synth2_19_), .Y(_4177_) );
	NOR2X1 NOR2X1_75 ( .A(_4133_), .B(_4177_), .Y(_4178_) );
	NOR2X1 NOR2X1_76 ( .A(micro_hash_synth_2_c_3_), .B(Hhash_synth2_19_), .Y(_4179_) );
	NOR2X1 NOR2X1_77 ( .A(_4179_), .B(_4178_), .Y(_4180_) );
	XOR2X1 XOR2X1_3 ( .A(_4176_), .B(_4180_), .Y(_4181_) );
	OAI21X1 OAI21X1_144 ( .A(Hhash_synth2_19_), .B(_3332__bF_buf2), .C(_3320_), .Y(_4182_) );
	OAI21X1 OAI21X1_145 ( .A(_3317_), .B(_4181_), .C(_4182_), .Y(_3047__19_) );
	XOR2X1 XOR2X1_4 ( .A(micro_hash_synth_2_c_4_), .B(Hhash_synth2_20_), .Y(_4183_) );
	INVX1 INVX1_63 ( .A(_4183_), .Y(_4184_) );
	OAI21X1 OAI21X1_146 ( .A(_4133_), .B(_4177_), .C(_4176_), .Y(_4185_) );
	OAI21X1 OAI21X1_147 ( .A(micro_hash_synth_2_c_3_), .B(Hhash_synth2_19_), .C(_4185_), .Y(_4186_) );
	NAND2X1 NAND2X1_126 ( .A(_4184_), .B(_4186_), .Y(_4187_) );
	NOR2X1 NOR2X1_78 ( .A(_4184_), .B(_4186_), .Y(_4188_) );
	INVX1 INVX1_64 ( .A(_4188_), .Y(_4189_) );
	NAND2X1 NAND2X1_127 ( .A(_4187_), .B(_4189_), .Y(_4190_) );
	OAI21X1 OAI21X1_148 ( .A(Hhash_synth2_20_), .B(_3332__bF_buf1), .C(_3320_), .Y(_4191_) );
	OAI21X1 OAI21X1_149 ( .A(_4190_), .B(_3317_), .C(_4191_), .Y(_3047__20_) );
	OAI21X1 OAI21X1_150 ( .A(Hhash_synth2_21_), .B(_3332__bF_buf0), .C(_3320_), .Y(_4192_) );
	AOI21X1 AOI21X1_70 ( .A(micro_hash_synth_2_c_4_), .B(Hhash_synth2_20_), .C(_4188_), .Y(_4193_) );
	INVX1 INVX1_65 ( .A(Hhash_synth2_21_), .Y(_4194_) );
	NOR2X1 NOR2X1_79 ( .A(_4144_), .B(_4194_), .Y(_4195_) );
	NOR2X1 NOR2X1_80 ( .A(micro_hash_synth_2_c_5_), .B(Hhash_synth2_21_), .Y(_4196_) );
	NOR2X1 NOR2X1_81 ( .A(_4196_), .B(_4195_), .Y(_4197_) );
	XOR2X1 XOR2X1_5 ( .A(_4193_), .B(_4197_), .Y(_4198_) );
	OAI21X1 OAI21X1_151 ( .A(_4198_), .B(_3317_), .C(_4192_), .Y(_3047__21_) );
	OAI21X1 OAI21X1_152 ( .A(Hhash_synth2_22_), .B(_3332__bF_buf3), .C(_3320_), .Y(_4199_) );
	XOR2X1 XOR2X1_6 ( .A(micro_hash_synth_2_c_6_), .B(Hhash_synth2_22_), .Y(_4200_) );
	INVX1 INVX1_66 ( .A(_4195_), .Y(_4201_) );
	OAI21X1 OAI21X1_153 ( .A(_4193_), .B(_4196_), .C(_4201_), .Y(_4202_) );
	NOR2X1 NOR2X1_82 ( .A(_4200_), .B(_4202_), .Y(_4203_) );
	NAND2X1 NAND2X1_128 ( .A(_4200_), .B(_4202_), .Y(_4204_) );
	NAND2X1 NAND2X1_129 ( .A(_3316__bF_buf0), .B(_4204_), .Y(_4205_) );
	OAI21X1 OAI21X1_154 ( .A(_4205_), .B(_4203_), .C(_4199_), .Y(_3047__22_) );
	OAI21X1 OAI21X1_155 ( .A(Hhash_synth2_23_), .B(_3332__bF_buf2), .C(_3320_), .Y(_4206_) );
	INVX1 INVX1_67 ( .A(Hhash_synth2_22_), .Y(_4207_) );
	OAI21X1 OAI21X1_156 ( .A(_4148_), .B(_4207_), .C(_4204_), .Y(_4208_) );
	XNOR2X1 XNOR2X1_6 ( .A(micro_hash_synth_2_c_7_), .B(Hhash_synth2_23_), .Y(_4209_) );
	INVX1 INVX1_68 ( .A(_4209_), .Y(_4210_) );
	AND2X2 AND2X2_30 ( .A(_4208_), .B(_4210_), .Y(_4211_) );
	OAI21X1 OAI21X1_157 ( .A(_4208_), .B(_4210_), .C(_3316__bF_buf3), .Y(_4212_) );
	OAI21X1 OAI21X1_158 ( .A(_4211_), .B(_4212_), .C(_4206_), .Y(_3047__23_) );
	NAND3X1 NAND3X1_53 ( .A(_3322_), .B(_3375_), .C(_3424__bF_buf2), .Y(_4213_) );
	OAI21X1 OAI21X1_159 ( .A(micro_hash_synth_2_x_0_), .B(_3424__bF_buf1), .C(_4213_), .Y(_4214_) );
	XNOR2X1 XNOR2X1_7 ( .A(micro_hash_synth_2_b_0_), .B(micro_hash_synth_2_a_0_), .Y(_4215_) );
	NAND2X1 NAND2X1_130 ( .A(_3432_), .B(_3333__bF_buf0), .Y(_4216_) );
	OAI22X1 OAI22X1_34 ( .A(_4215_), .B(_4216_), .C(_4214_), .D(_3437_), .Y(_3053__0_) );
	NAND3X1 NAND3X1_54 ( .A(_3325_), .B(_3378_), .C(_3424__bF_buf0), .Y(_4217_) );
	OAI21X1 OAI21X1_160 ( .A(micro_hash_synth_2_x_1_), .B(_3424__bF_buf3), .C(_4217_), .Y(_4218_) );
	XNOR2X1 XNOR2X1_8 ( .A(micro_hash_synth_2_b_1_), .B(micro_hash_synth_2_a_1_), .Y(_4219_) );
	OAI22X1 OAI22X1_35 ( .A(_4216_), .B(_4219_), .C(_4218_), .D(_3437_), .Y(_3053__1_) );
	NAND3X1 NAND3X1_55 ( .A(_4115_), .B(_4128_), .C(_3424__bF_buf2), .Y(_4220_) );
	OAI21X1 OAI21X1_161 ( .A(micro_hash_synth_2_x_2_), .B(_3424__bF_buf1), .C(_4220_), .Y(_4221_) );
	XNOR2X1 XNOR2X1_9 ( .A(micro_hash_synth_2_b_2_), .B(micro_hash_synth_2_a_2_), .Y(_4222_) );
	OAI22X1 OAI22X1_36 ( .A(_4216_), .B(_4222_), .C(_4221_), .D(_3437_), .Y(_3053__2_) );
	XOR2X1 XOR2X1_7 ( .A(micro_hash_synth_2_b_3_), .B(micro_hash_synth_2_a_3_), .Y(_4223_) );
	OAI21X1 OAI21X1_162 ( .A(_3332__bF_buf1), .B(_4223_), .C(_3437_), .Y(_4224_) );
	OAI21X1 OAI21X1_163 ( .A(micro_hash_synth_2_b_3_), .B(micro_hash_synth_2_a_3_), .C(_3424__bF_buf0), .Y(_4225_) );
	OAI21X1 OAI21X1_164 ( .A(_3719_), .B(_3424__bF_buf3), .C(_4225_), .Y(_4226_) );
	NAND2X1 NAND2X1_131 ( .A(_3431_), .B(_4226_), .Y(_4227_) );
	NAND2X1 NAND2X1_132 ( .A(_4224_), .B(_4227_), .Y(_3053__3_) );
	NAND3X1 NAND3X1_56 ( .A(_4140_), .B(_4137_), .C(_3424__bF_buf2), .Y(_4228_) );
	OAI21X1 OAI21X1_165 ( .A(micro_hash_synth_2_x_4_), .B(_3424__bF_buf1), .C(_4228_), .Y(_4229_) );
	XNOR2X1 XNOR2X1_10 ( .A(micro_hash_synth_2_b_4_), .B(micro_hash_synth_2_a_4_), .Y(_4230_) );
	OAI22X1 OAI22X1_37 ( .A(_4216_), .B(_4230_), .C(_4229_), .D(_3437_), .Y(_3053__4_) );
	NOR2X1 NOR2X1_83 ( .A(micro_hash_synth_2_b_5_), .B(micro_hash_synth_2_a_5_), .Y(_4231_) );
	OAI21X1 OAI21X1_166 ( .A(_3311_), .B(_3313_), .C(_4231_), .Y(_4232_) );
	OAI21X1 OAI21X1_167 ( .A(micro_hash_synth_2_x_5_), .B(_3424__bF_buf0), .C(_4232_), .Y(_4233_) );
	XNOR2X1 XNOR2X1_11 ( .A(micro_hash_synth_2_b_5_), .B(micro_hash_synth_2_a_5_), .Y(_4234_) );
	OAI22X1 OAI22X1_38 ( .A(_4216_), .B(_4234_), .C(_4233_), .D(_3437_), .Y(_3053__5_) );
	NOR2X1 NOR2X1_84 ( .A(micro_hash_synth_2_b_6_), .B(micro_hash_synth_2_a_6_), .Y(_4235_) );
	OAI21X1 OAI21X1_168 ( .A(_3311_), .B(_3313_), .C(_4235_), .Y(_4236_) );
	OAI21X1 OAI21X1_169 ( .A(micro_hash_synth_2_x_6_), .B(_3424__bF_buf3), .C(_4236_), .Y(_4237_) );
	XNOR2X1 XNOR2X1_12 ( .A(micro_hash_synth_2_b_6_), .B(micro_hash_synth_2_a_6_), .Y(_4238_) );
	OAI22X1 OAI22X1_39 ( .A(_4216_), .B(_4238_), .C(_4237_), .D(_3437_), .Y(_3053__6_) );
	XOR2X1 XOR2X1_8 ( .A(micro_hash_synth_2_b_7_), .B(micro_hash_synth_2_a_7_), .Y(_4239_) );
	OAI21X1 OAI21X1_170 ( .A(_3332__bF_buf0), .B(_4239_), .C(_3437_), .Y(_4240_) );
	NAND2X1 NAND2X1_133 ( .A(_4121_), .B(_4152_), .Y(_4241_) );
	NOR2X1 NOR2X1_85 ( .A(_4241_), .B(_3436_), .Y(_4242_) );
	OAI21X1 OAI21X1_171 ( .A(_3424__bF_buf2), .B(micro_hash_synth_2_x_7_), .C(_3431_), .Y(_4243_) );
	OAI21X1 OAI21X1_172 ( .A(_4243_), .B(_4242_), .C(_4240_), .Y(_3053__7_) );
	INVX1 INVX1_69 ( .A(micro_hash_synth_2_W_24__0_), .Y(_4244_) );
	XOR2X1 XOR2X1_9 ( .A(micro_hash_synth_2_W_10__0_), .B(micro_hash_synth_2_W_15__0_), .Y(_4245_) );
	NOR2X1 NOR2X1_86 ( .A(micro_hash_synth_2_W_21__0_), .B(_4245_), .Y(_4246_) );
	OAI22X1 OAI22X1_40 ( .A(_4735__bF_buf15), .B(_4246_), .C(_4740__bF_buf13), .D(_4244_), .Y(_3216_) );
	INVX1 INVX1_70 ( .A(micro_hash_synth_2_W_21__1_), .Y(_4247_) );
	OAI21X1 OAI21X1_173 ( .A(_3546_), .B(micro_hash_synth_2_W_15__1_), .C(_4247_), .Y(_4248_) );
	AOI21X1 AOI21X1_71 ( .A(_3546_), .B(micro_hash_synth_2_W_15__1_), .C(_4248_), .Y(_4249_) );
	OAI22X1 OAI22X1_41 ( .A(_4735__bF_buf14), .B(_4249_), .C(_4740__bF_buf12), .D(_3533_), .Y(_3217_) );
	INVX1 INVX1_71 ( .A(micro_hash_synth_2_W_21__2_), .Y(_4250_) );
	OAI21X1 OAI21X1_174 ( .A(_3646_), .B(micro_hash_synth_2_W_15__2_), .C(_4250_), .Y(_4251_) );
	AOI21X1 AOI21X1_72 ( .A(_3646_), .B(micro_hash_synth_2_W_15__2_), .C(_4251_), .Y(_4252_) );
	OAI22X1 OAI22X1_42 ( .A(_4735__bF_buf13), .B(_4252_), .C(_4740__bF_buf11), .D(_3629_), .Y(_3218_) );
	INVX1 INVX1_72 ( .A(micro_hash_synth_2_W_21__3_), .Y(_4253_) );
	OAI21X1 OAI21X1_175 ( .A(_3761_), .B(micro_hash_synth_2_W_15__3_), .C(_4253_), .Y(_4254_) );
	AOI21X1 AOI21X1_73 ( .A(_3761_), .B(micro_hash_synth_2_W_15__3_), .C(_4254_), .Y(_4255_) );
	OAI22X1 OAI22X1_43 ( .A(_4735__bF_buf12), .B(_4255_), .C(_4740__bF_buf10), .D(_3729_), .Y(_3219_) );
	INVX1 INVX1_73 ( .A(micro_hash_synth_2_W_21__4_), .Y(_4256_) );
	OAI21X1 OAI21X1_176 ( .A(_3827_), .B(micro_hash_synth_2_W_15__4_), .C(_4256_), .Y(_4257_) );
	AOI21X1 AOI21X1_74 ( .A(_3827_), .B(micro_hash_synth_2_W_15__4_), .C(_4257_), .Y(_4258_) );
	OAI22X1 OAI22X1_44 ( .A(_4735__bF_buf11), .B(_4258_), .C(_4740__bF_buf9), .D(_3813_), .Y(_3220_) );
	INVX1 INVX1_74 ( .A(micro_hash_synth_2_W_21__5_), .Y(_4259_) );
	OAI21X1 OAI21X1_177 ( .A(_3929_), .B(micro_hash_synth_2_W_15__5_), .C(_4259_), .Y(_4260_) );
	AOI21X1 AOI21X1_75 ( .A(_3929_), .B(micro_hash_synth_2_W_15__5_), .C(_4260_), .Y(_4261_) );
	OAI22X1 OAI22X1_45 ( .A(_4735__bF_buf10), .B(_4261_), .C(_4740__bF_buf8), .D(_3915_), .Y(_3221_) );
	INVX1 INVX1_75 ( .A(micro_hash_synth_2_W_21__6_), .Y(_4262_) );
	OAI21X1 OAI21X1_178 ( .A(_4015_), .B(micro_hash_synth_2_W_15__6_), .C(_4262_), .Y(_4263_) );
	AOI21X1 AOI21X1_76 ( .A(_4015_), .B(micro_hash_synth_2_W_15__6_), .C(_4263_), .Y(_4264_) );
	OAI22X1 OAI22X1_46 ( .A(_4735__bF_buf9), .B(_4264_), .C(_4740__bF_buf7), .D(_3996_), .Y(_3223_) );
	INVX1 INVX1_76 ( .A(micro_hash_synth_2_W_10__7_), .Y(_4265_) );
	INVX1 INVX1_77 ( .A(micro_hash_synth_2_W_21__7_), .Y(_4266_) );
	OAI21X1 OAI21X1_179 ( .A(_4265_), .B(micro_hash_synth_2_W_15__7_), .C(_4266_), .Y(_4267_) );
	AOI21X1 AOI21X1_77 ( .A(_4265_), .B(micro_hash_synth_2_W_15__7_), .C(_4267_), .Y(_4268_) );
	OAI22X1 OAI22X1_47 ( .A(_4735__bF_buf8), .B(_4268_), .C(_4740__bF_buf6), .D(_4068_), .Y(_3224_) );
	INVX8 INVX8_1 ( .A(_4740__bF_buf5), .Y(_4269_) );
	NAND2X1 NAND2X1_134 ( .A(micro_hash_synth_2_W_23__0_), .B(_4269__bF_buf6), .Y(_4270_) );
	XOR2X1 XOR2X1_10 ( .A(micro_hash_synth_2_W_9__0_), .B(micro_hash_synth_2_W_14__0_), .Y(_4271_) );
	NOR2X1 NOR2X1_87 ( .A(micro_hash_synth_2_W_20__0_), .B(_4271_), .Y(_4272_) );
	OAI21X1 OAI21X1_180 ( .A(_4735__bF_buf7), .B(_4272_), .C(_4270_), .Y(_3225_) );
	XOR2X1 XOR2X1_11 ( .A(micro_hash_synth_2_W_9__1_), .B(micro_hash_synth_2_W_14__1_), .Y(_4273_) );
	NOR2X1 NOR2X1_88 ( .A(micro_hash_synth_2_W_20__1_), .B(_4273_), .Y(_4274_) );
	OAI22X1 OAI22X1_48 ( .A(_4735__bF_buf6), .B(_4274_), .C(_4740__bF_buf4), .D(_4745_), .Y(_3226_) );
	XOR2X1 XOR2X1_12 ( .A(micro_hash_synth_2_W_9__2_), .B(micro_hash_synth_2_W_14__2_), .Y(_4275_) );
	NOR2X1 NOR2X1_89 ( .A(micro_hash_synth_2_W_20__2_), .B(_4275_), .Y(_4276_) );
	OAI22X1 OAI22X1_49 ( .A(_4735__bF_buf5), .B(_4276_), .C(_4740__bF_buf3), .D(_4750_), .Y(_3227_) );
	NAND2X1 NAND2X1_135 ( .A(micro_hash_synth_2_W_23__3_), .B(_4269__bF_buf5), .Y(_4277_) );
	XOR2X1 XOR2X1_13 ( .A(micro_hash_synth_2_W_9__3_), .B(micro_hash_synth_2_W_14__3_), .Y(_4278_) );
	NOR2X1 NOR2X1_90 ( .A(micro_hash_synth_2_W_20__3_), .B(_4278_), .Y(_4279_) );
	OAI21X1 OAI21X1_181 ( .A(_4735__bF_buf4), .B(_4279_), .C(_4277_), .Y(_3228_) );
	NAND2X1 NAND2X1_136 ( .A(micro_hash_synth_2_W_23__4_), .B(_4269__bF_buf4), .Y(_4280_) );
	XOR2X1 XOR2X1_14 ( .A(micro_hash_synth_2_W_9__4_), .B(micro_hash_synth_2_W_14__4_), .Y(_4281_) );
	NOR2X1 NOR2X1_91 ( .A(micro_hash_synth_2_W_20__4_), .B(_4281_), .Y(_4282_) );
	OAI21X1 OAI21X1_182 ( .A(_4735__bF_buf3), .B(_4282_), .C(_4280_), .Y(_3229_) );
	NAND2X1 NAND2X1_137 ( .A(micro_hash_synth_2_W_23__5_), .B(_4269__bF_buf3), .Y(_4283_) );
	XOR2X1 XOR2X1_15 ( .A(micro_hash_synth_2_W_9__5_), .B(micro_hash_synth_2_W_14__5_), .Y(_4284_) );
	NOR2X1 NOR2X1_92 ( .A(micro_hash_synth_2_W_20__5_), .B(_4284_), .Y(_4285_) );
	OAI21X1 OAI21X1_183 ( .A(_4735__bF_buf2), .B(_4285_), .C(_4283_), .Y(_3230_) );
	INVX1 INVX1_78 ( .A(micro_hash_synth_2_W_20__6_), .Y(_4286_) );
	OAI21X1 OAI21X1_184 ( .A(_4012_), .B(micro_hash_synth_2_W_14__6_), .C(_4286_), .Y(_4287_) );
	AOI21X1 AOI21X1_78 ( .A(_4012_), .B(micro_hash_synth_2_W_14__6_), .C(_4287_), .Y(_4288_) );
	OAI22X1 OAI22X1_50 ( .A(_4735__bF_buf1), .B(_4288_), .C(_4740__bF_buf2), .D(_4764_), .Y(_3231_) );
	XOR2X1 XOR2X1_16 ( .A(micro_hash_synth_2_W_9__7_), .B(micro_hash_synth_2_W_14__7_), .Y(_4289_) );
	NOR2X1 NOR2X1_93 ( .A(micro_hash_synth_2_W_20__7_), .B(_4289_), .Y(_4290_) );
	OAI22X1 OAI22X1_51 ( .A(_4735__bF_buf0), .B(_4290_), .C(_4740__bF_buf1), .D(_4769_), .Y(_3232_) );
	INVX1 INVX1_79 ( .A(micro_hash_synth_2_W_7__0_), .Y(_4291_) );
	INVX1 INVX1_80 ( .A(bloque_in_1_56_), .Y(_4292_) );
	OAI22X1 OAI22X1_52 ( .A(_4292_), .B(_4735__bF_buf15), .C(_4740__bF_buf0), .D(_4291_), .Y(_3234_) );
	INVX1 INVX1_81 ( .A(bloque_in_1_57_), .Y(_4293_) );
	OAI22X1 OAI22X1_53 ( .A(_4293_), .B(_4735__bF_buf14), .C(_4740__bF_buf13), .D(_3560_), .Y(_3235_) );
	INVX1 INVX1_82 ( .A(bloque_in_1_58_), .Y(_4294_) );
	OAI22X1 OAI22X1_54 ( .A(_4294_), .B(_4735__bF_buf13), .C(_4740__bF_buf12), .D(_3694_), .Y(_3236_) );
	INVX1 INVX1_83 ( .A(micro_hash_synth_2_W_7__3_), .Y(_4295_) );
	INVX1 INVX1_84 ( .A(bloque_in_1_59_), .Y(_4296_) );
	OAI22X1 OAI22X1_55 ( .A(_4296_), .B(_4735__bF_buf12), .C(_4740__bF_buf11), .D(_4295_), .Y(_3237_) );
	INVX1 INVX1_85 ( .A(micro_hash_synth_2_W_7__4_), .Y(_4297_) );
	INVX1 INVX1_86 ( .A(bloque_in_1_60_), .Y(_4298_) );
	OAI22X1 OAI22X1_56 ( .A(_4298_), .B(_4735__bF_buf11), .C(_4740__bF_buf10), .D(_4297_), .Y(_3238_) );
	INVX1 INVX1_87 ( .A(micro_hash_synth_2_W_7__5_), .Y(_4299_) );
	INVX1 INVX1_88 ( .A(bloque_in_1_61_), .Y(_4300_) );
	OAI22X1 OAI22X1_57 ( .A(_4300_), .B(_4735__bF_buf10), .C(_4740__bF_buf9), .D(_4299_), .Y(_3239_) );
	INVX1 INVX1_89 ( .A(bloque_in_1_62_), .Y(_4301_) );
	OAI22X1 OAI22X1_58 ( .A(_4301_), .B(_4735__bF_buf9), .C(_4740__bF_buf8), .D(_4022_), .Y(_3240_) );
	INVX1 INVX1_90 ( .A(micro_hash_synth_2_W_7__7_), .Y(_4302_) );
	INVX1 INVX1_91 ( .A(bloque_in_1_63_), .Y(_4303_) );
	OAI22X1 OAI22X1_59 ( .A(_4303_), .B(_4735__bF_buf8), .C(_4740__bF_buf7), .D(_4302_), .Y(_3241_) );
	NAND2X1 NAND2X1_138 ( .A(micro_hash_synth_2_W_22__0_), .B(_4269__bF_buf2), .Y(_4304_) );
	INVX1 INVX1_92 ( .A(micro_hash_synth_2_W_19__0_), .Y(_4305_) );
	OAI21X1 OAI21X1_185 ( .A(_4800_), .B(micro_hash_synth_2_W_13__0_), .C(_4305_), .Y(_4306_) );
	AOI21X1 AOI21X1_79 ( .A(_4800_), .B(micro_hash_synth_2_W_13__0_), .C(_4306_), .Y(_4307_) );
	OAI21X1 OAI21X1_186 ( .A(_4735__bF_buf7), .B(_4307_), .C(_4304_), .Y(_3242_) );
	INVX1 INVX1_93 ( .A(micro_hash_synth_2_W_19__1_), .Y(_4308_) );
	OAI21X1 OAI21X1_187 ( .A(_4802_), .B(micro_hash_synth_2_W_13__1_), .C(_4308_), .Y(_4309_) );
	AOI21X1 AOI21X1_80 ( .A(_4802_), .B(micro_hash_synth_2_W_13__1_), .C(_4309_), .Y(_4310_) );
	OAI22X1 OAI22X1_60 ( .A(_4735__bF_buf6), .B(_4310_), .C(_4740__bF_buf6), .D(_4777_), .Y(_3243_) );
	INVX1 INVX1_94 ( .A(micro_hash_synth_2_W_19__2_), .Y(_4311_) );
	OAI21X1 OAI21X1_188 ( .A(_4804_), .B(micro_hash_synth_2_W_13__2_), .C(_4311_), .Y(_4312_) );
	AOI21X1 AOI21X1_81 ( .A(_4804_), .B(micro_hash_synth_2_W_13__2_), .C(_4312_), .Y(_4313_) );
	OAI22X1 OAI22X1_61 ( .A(_4735__bF_buf5), .B(_4313_), .C(_4740__bF_buf5), .D(_4782_), .Y(_3245_) );
	NAND2X1 NAND2X1_139 ( .A(micro_hash_synth_2_W_22__3_), .B(_4269__bF_buf1), .Y(_4314_) );
	INVX1 INVX1_95 ( .A(micro_hash_synth_2_W_19__3_), .Y(_4315_) );
	OAI21X1 OAI21X1_189 ( .A(_4806_), .B(micro_hash_synth_2_W_13__3_), .C(_4315_), .Y(_4316_) );
	AOI21X1 AOI21X1_82 ( .A(_4806_), .B(micro_hash_synth_2_W_13__3_), .C(_4316_), .Y(_4317_) );
	OAI21X1 OAI21X1_190 ( .A(_4735__bF_buf4), .B(_4317_), .C(_4314_), .Y(_3246_) );
	NAND2X1 NAND2X1_140 ( .A(micro_hash_synth_2_W_22__4_), .B(_4269__bF_buf0), .Y(_4318_) );
	INVX1 INVX1_96 ( .A(micro_hash_synth_2_W_19__4_), .Y(_4319_) );
	OAI21X1 OAI21X1_191 ( .A(_4808_), .B(micro_hash_synth_2_W_13__4_), .C(_4319_), .Y(_4320_) );
	AOI21X1 AOI21X1_83 ( .A(_4808_), .B(micro_hash_synth_2_W_13__4_), .C(_4320_), .Y(_4321_) );
	OAI21X1 OAI21X1_192 ( .A(_4735__bF_buf3), .B(_4321_), .C(_4318_), .Y(_3247_) );
	NAND2X1 NAND2X1_141 ( .A(micro_hash_synth_2_W_22__5_), .B(_4269__bF_buf6), .Y(_4322_) );
	INVX1 INVX1_97 ( .A(micro_hash_synth_2_W_19__5_), .Y(_4323_) );
	OAI21X1 OAI21X1_193 ( .A(_4810_), .B(micro_hash_synth_2_W_13__5_), .C(_4323_), .Y(_4324_) );
	AOI21X1 AOI21X1_84 ( .A(_4810_), .B(micro_hash_synth_2_W_13__5_), .C(_4324_), .Y(_4325_) );
	OAI21X1 OAI21X1_194 ( .A(_4735__bF_buf2), .B(_4325_), .C(_4322_), .Y(_3248_) );
	NAND2X1 NAND2X1_142 ( .A(micro_hash_synth_2_W_22__6_), .B(_4269__bF_buf5), .Y(_4326_) );
	INVX1 INVX1_98 ( .A(micro_hash_synth_2_W_19__6_), .Y(_4327_) );
	OAI21X1 OAI21X1_195 ( .A(_4812_), .B(micro_hash_synth_2_W_13__6_), .C(_4327_), .Y(_4328_) );
	AOI21X1 AOI21X1_85 ( .A(_4812_), .B(micro_hash_synth_2_W_13__6_), .C(_4328_), .Y(_4329_) );
	OAI21X1 OAI21X1_196 ( .A(_4735__bF_buf1), .B(_4329_), .C(_4326_), .Y(_3249_) );
	NAND2X1 NAND2X1_143 ( .A(micro_hash_synth_2_W_22__7_), .B(_4269__bF_buf4), .Y(_4330_) );
	INVX1 INVX1_99 ( .A(micro_hash_synth_2_W_19__7_), .Y(_4331_) );
	OAI21X1 OAI21X1_197 ( .A(_4814_), .B(micro_hash_synth_2_W_13__7_), .C(_4331_), .Y(_4332_) );
	AOI21X1 AOI21X1_86 ( .A(_4814_), .B(micro_hash_synth_2_W_13__7_), .C(_4332_), .Y(_4333_) );
	OAI21X1 OAI21X1_198 ( .A(_4735__bF_buf0), .B(_4333_), .C(_4330_), .Y(_3250_) );
	INVX1 INVX1_100 ( .A(bloque_in_1_72_), .Y(_4334_) );
	NAND2X1 NAND2X1_144 ( .A(micro_hash_synth_2_W_9__0_), .B(_4269__bF_buf3), .Y(_4335_) );
	OAI21X1 OAI21X1_199 ( .A(_4334_), .B(_4735__bF_buf15), .C(_4335_), .Y(_3251_) );
	INVX1 INVX1_101 ( .A(bloque_in_1_73_), .Y(_4336_) );
	NAND2X1 NAND2X1_145 ( .A(micro_hash_synth_2_W_9__1_), .B(_4269__bF_buf2), .Y(_4337_) );
	OAI21X1 OAI21X1_200 ( .A(_4336_), .B(_4735__bF_buf14), .C(_4337_), .Y(_3252_) );
	INVX1 INVX1_102 ( .A(bloque_in_1_74_), .Y(_4338_) );
	NAND2X1 NAND2X1_146 ( .A(micro_hash_synth_2_W_9__2_), .B(_4269__bF_buf1), .Y(_4339_) );
	OAI21X1 OAI21X1_201 ( .A(_4338_), .B(_4735__bF_buf13), .C(_4339_), .Y(_3253_) );
	INVX1 INVX1_103 ( .A(bloque_in_1_75_), .Y(_4340_) );
	NAND2X1 NAND2X1_147 ( .A(micro_hash_synth_2_W_9__3_), .B(_4269__bF_buf0), .Y(_4341_) );
	OAI21X1 OAI21X1_202 ( .A(_4340_), .B(_4735__bF_buf12), .C(_4341_), .Y(_3254_) );
	INVX1 INVX1_104 ( .A(bloque_in_1_76_), .Y(_4342_) );
	NAND2X1 NAND2X1_148 ( .A(micro_hash_synth_2_W_9__4_), .B(_4269__bF_buf6), .Y(_4343_) );
	OAI21X1 OAI21X1_203 ( .A(_4342_), .B(_4735__bF_buf11), .C(_4343_), .Y(_3256_) );
	INVX1 INVX1_105 ( .A(bloque_in_1_77_), .Y(_4344_) );
	NAND2X1 NAND2X1_149 ( .A(micro_hash_synth_2_W_9__5_), .B(_4269__bF_buf5), .Y(_4345_) );
	OAI21X1 OAI21X1_204 ( .A(_4344_), .B(_4735__bF_buf10), .C(_4345_), .Y(_3257_) );
	INVX1 INVX1_106 ( .A(bloque_in_1_78_), .Y(_4346_) );
	OAI22X1 OAI22X1_62 ( .A(_4346_), .B(_4735__bF_buf9), .C(_4740__bF_buf4), .D(_4012_), .Y(_3258_) );
	INVX1 INVX1_107 ( .A(bloque_in_1_79_), .Y(_4347_) );
	NAND2X1 NAND2X1_150 ( .A(micro_hash_synth_2_W_9__7_), .B(_4269__bF_buf4), .Y(_4348_) );
	OAI21X1 OAI21X1_205 ( .A(_4347_), .B(_4735__bF_buf8), .C(_4348_), .Y(_3259_) );
	INVX1 INVX1_108 ( .A(micro_hash_synth_2_W_4__0_), .Y(_4349_) );
	INVX1 INVX1_109 ( .A(bloque_in_1_32_), .Y(_4350_) );
	OAI22X1 OAI22X1_63 ( .A(_4350_), .B(_4735__bF_buf7), .C(_4740__bF_buf3), .D(_4349_), .Y(_3260_) );
	INVX1 INVX1_110 ( .A(micro_hash_synth_2_W_4__1_), .Y(_4351_) );
	INVX1 INVX1_111 ( .A(bloque_in_1_33_), .Y(_4352_) );
	OAI22X1 OAI22X1_64 ( .A(_4352_), .B(_4735__bF_buf6), .C(_4740__bF_buf2), .D(_4351_), .Y(_3261_) );
	INVX1 INVX1_112 ( .A(micro_hash_synth_2_W_4__2_), .Y(_4353_) );
	INVX1 INVX1_113 ( .A(bloque_in_1_34_), .Y(_4354_) );
	OAI22X1 OAI22X1_65 ( .A(_4354_), .B(_4735__bF_buf5), .C(_4740__bF_buf1), .D(_4353_), .Y(_3262_) );
	INVX1 INVX1_114 ( .A(micro_hash_synth_2_W_4__3_), .Y(_4355_) );
	INVX1 INVX1_115 ( .A(bloque_in_1_35_), .Y(_4356_) );
	OAI22X1 OAI22X1_66 ( .A(_4356_), .B(_4735__bF_buf4), .C(_4740__bF_buf0), .D(_4355_), .Y(_3263_) );
	INVX1 INVX1_116 ( .A(micro_hash_synth_2_W_4__4_), .Y(_4357_) );
	INVX1 INVX1_117 ( .A(bloque_in_1_36_), .Y(_4358_) );
	OAI22X1 OAI22X1_67 ( .A(_4358_), .B(_4735__bF_buf3), .C(_4740__bF_buf13), .D(_4357_), .Y(_3264_) );
	INVX1 INVX1_118 ( .A(micro_hash_synth_2_W_4__5_), .Y(_4359_) );
	INVX1 INVX1_119 ( .A(bloque_in_1_37_), .Y(_4360_) );
	OAI22X1 OAI22X1_68 ( .A(_4360_), .B(_4735__bF_buf2), .C(_4740__bF_buf12), .D(_4359_), .Y(_3265_) );
	INVX1 INVX1_120 ( .A(micro_hash_synth_2_W_4__6_), .Y(_4361_) );
	INVX1 INVX1_121 ( .A(bloque_in_1_38_), .Y(_4362_) );
	OAI22X1 OAI22X1_69 ( .A(_4362_), .B(_4735__bF_buf1), .C(_4740__bF_buf11), .D(_4361_), .Y(_3267_) );
	INVX1 INVX1_122 ( .A(micro_hash_synth_2_W_4__7_), .Y(_4363_) );
	INVX1 INVX1_123 ( .A(bloque_in_1_39_), .Y(_4364_) );
	OAI22X1 OAI22X1_70 ( .A(_4364_), .B(_4735__bF_buf0), .C(_4740__bF_buf10), .D(_4363_), .Y(_3268_) );
	NAND2X1 NAND2X1_151 ( .A(micro_hash_synth_2_W_21__0_), .B(_4269__bF_buf3), .Y(_4365_) );
	OAI21X1 OAI21X1_206 ( .A(_4291_), .B(micro_hash_synth_2_W_12__0_), .C(_3480_), .Y(_4366_) );
	AOI21X1 AOI21X1_87 ( .A(micro_hash_synth_2_W_12__0_), .B(_4291_), .C(_4366_), .Y(_4367_) );
	OAI21X1 OAI21X1_207 ( .A(_4735__bF_buf15), .B(_4367_), .C(_4365_), .Y(_3269_) );
	OAI21X1 OAI21X1_208 ( .A(_3560_), .B(micro_hash_synth_2_W_12__1_), .C(_3513_), .Y(_4368_) );
	AOI21X1 AOI21X1_88 ( .A(micro_hash_synth_2_W_12__1_), .B(_3560_), .C(_4368_), .Y(_4369_) );
	OAI22X1 OAI22X1_71 ( .A(_4735__bF_buf14), .B(_4369_), .C(_4740__bF_buf9), .D(_4247_), .Y(_3270_) );
	OAI21X1 OAI21X1_209 ( .A(_3694_), .B(micro_hash_synth_2_W_12__2_), .C(_3614_), .Y(_4370_) );
	AOI21X1 AOI21X1_89 ( .A(micro_hash_synth_2_W_12__2_), .B(_3694_), .C(_4370_), .Y(_4371_) );
	OAI22X1 OAI22X1_72 ( .A(_4735__bF_buf13), .B(_4371_), .C(_4740__bF_buf8), .D(_4250_), .Y(_3271_) );
	OAI21X1 OAI21X1_210 ( .A(_4295_), .B(micro_hash_synth_2_W_12__3_), .C(_3744_), .Y(_4372_) );
	AOI21X1 AOI21X1_90 ( .A(micro_hash_synth_2_W_12__3_), .B(_4295_), .C(_4372_), .Y(_4373_) );
	OAI22X1 OAI22X1_73 ( .A(_4735__bF_buf12), .B(_4373_), .C(_4740__bF_buf7), .D(_4253_), .Y(_3272_) );
	OAI21X1 OAI21X1_211 ( .A(_4297_), .B(micro_hash_synth_2_W_12__4_), .C(_3841_), .Y(_4374_) );
	AOI21X1 AOI21X1_91 ( .A(micro_hash_synth_2_W_12__4_), .B(_4297_), .C(_4374_), .Y(_4375_) );
	OAI22X1 OAI22X1_74 ( .A(_4735__bF_buf11), .B(_4375_), .C(_4740__bF_buf6), .D(_4256_), .Y(_3273_) );
	OAI21X1 OAI21X1_212 ( .A(_4299_), .B(micro_hash_synth_2_W_12__5_), .C(_3898_), .Y(_4376_) );
	AOI21X1 AOI21X1_92 ( .A(micro_hash_synth_2_W_12__5_), .B(_4299_), .C(_4376_), .Y(_4377_) );
	OAI22X1 OAI22X1_75 ( .A(_4735__bF_buf10), .B(_4377_), .C(_4740__bF_buf5), .D(_4259_), .Y(_3274_) );
	OAI21X1 OAI21X1_213 ( .A(_4022_), .B(micro_hash_synth_2_W_12__6_), .C(_3982_), .Y(_4378_) );
	AOI21X1 AOI21X1_93 ( .A(micro_hash_synth_2_W_12__6_), .B(_4022_), .C(_4378_), .Y(_4379_) );
	OAI22X1 OAI22X1_76 ( .A(_4735__bF_buf9), .B(_4379_), .C(_4740__bF_buf4), .D(_4262_), .Y(_3275_) );
	OAI21X1 OAI21X1_214 ( .A(_4302_), .B(micro_hash_synth_2_W_12__7_), .C(_4052_), .Y(_4380_) );
	AOI21X1 AOI21X1_94 ( .A(micro_hash_synth_2_W_12__7_), .B(_4302_), .C(_4380_), .Y(_4381_) );
	OAI22X1 OAI22X1_77 ( .A(_4735__bF_buf8), .B(_4381_), .C(_4740__bF_buf3), .D(_4266_), .Y(_3276_) );
	NAND2X1 NAND2X1_152 ( .A(micro_hash_synth_2_W_20__0_), .B(_4269__bF_buf2), .Y(_4382_) );
	INVX1 INVX1_124 ( .A(micro_hash_synth_2_W_6__0_), .Y(_4383_) );
	INVX1 INVX1_125 ( .A(micro_hash_synth_2_W_17__0_), .Y(_4384_) );
	OAI21X1 OAI21X1_215 ( .A(_4383_), .B(micro_hash_synth_2_W_11__0_), .C(_4384_), .Y(_4385_) );
	AOI21X1 AOI21X1_95 ( .A(micro_hash_synth_2_W_11__0_), .B(_4383_), .C(_4385_), .Y(_4386_) );
	OAI21X1 OAI21X1_216 ( .A(_4735__bF_buf7), .B(_4386_), .C(_4382_), .Y(_3278_) );
	NAND2X1 NAND2X1_153 ( .A(micro_hash_synth_2_W_20__1_), .B(_4269__bF_buf1), .Y(_4387_) );
	INVX1 INVX1_126 ( .A(micro_hash_synth_2_W_6__1_), .Y(_4388_) );
	INVX1 INVX1_127 ( .A(micro_hash_synth_2_W_17__1_), .Y(_4389_) );
	OAI21X1 OAI21X1_217 ( .A(_4388_), .B(micro_hash_synth_2_W_11__1_), .C(_4389_), .Y(_4390_) );
	AOI21X1 AOI21X1_96 ( .A(micro_hash_synth_2_W_11__1_), .B(_4388_), .C(_4390_), .Y(_4391_) );
	OAI21X1 OAI21X1_218 ( .A(_4735__bF_buf6), .B(_4391_), .C(_4387_), .Y(_3279_) );
	NAND2X1 NAND2X1_154 ( .A(micro_hash_synth_2_W_20__2_), .B(_4269__bF_buf0), .Y(_4392_) );
	INVX1 INVX1_128 ( .A(micro_hash_synth_2_W_6__2_), .Y(_4393_) );
	INVX1 INVX1_129 ( .A(micro_hash_synth_2_W_17__2_), .Y(_4394_) );
	OAI21X1 OAI21X1_219 ( .A(_4393_), .B(micro_hash_synth_2_W_11__2_), .C(_4394_), .Y(_4395_) );
	AOI21X1 AOI21X1_97 ( .A(micro_hash_synth_2_W_11__2_), .B(_4393_), .C(_4395_), .Y(_4396_) );
	OAI21X1 OAI21X1_220 ( .A(_4735__bF_buf5), .B(_4396_), .C(_4392_), .Y(_3280_) );
	NAND2X1 NAND2X1_155 ( .A(micro_hash_synth_2_W_20__3_), .B(_4269__bF_buf6), .Y(_4397_) );
	INVX1 INVX1_130 ( .A(micro_hash_synth_2_W_6__3_), .Y(_4398_) );
	INVX1 INVX1_131 ( .A(micro_hash_synth_2_W_17__3_), .Y(_4399_) );
	OAI21X1 OAI21X1_221 ( .A(_4398_), .B(micro_hash_synth_2_W_11__3_), .C(_4399_), .Y(_4400_) );
	AOI21X1 AOI21X1_98 ( .A(micro_hash_synth_2_W_11__3_), .B(_4398_), .C(_4400_), .Y(_4401_) );
	OAI21X1 OAI21X1_222 ( .A(_4735__bF_buf4), .B(_4401_), .C(_4397_), .Y(_3281_) );
	NAND2X1 NAND2X1_156 ( .A(micro_hash_synth_2_W_20__4_), .B(_4269__bF_buf5), .Y(_4402_) );
	INVX1 INVX1_132 ( .A(micro_hash_synth_2_W_6__4_), .Y(_4403_) );
	INVX1 INVX1_133 ( .A(micro_hash_synth_2_W_17__4_), .Y(_4404_) );
	OAI21X1 OAI21X1_223 ( .A(_4403_), .B(micro_hash_synth_2_W_11__4_), .C(_4404_), .Y(_4405_) );
	AOI21X1 AOI21X1_99 ( .A(micro_hash_synth_2_W_11__4_), .B(_4403_), .C(_4405_), .Y(_4406_) );
	OAI21X1 OAI21X1_224 ( .A(_4735__bF_buf3), .B(_4406_), .C(_4402_), .Y(_3282_) );
	NAND2X1 NAND2X1_157 ( .A(micro_hash_synth_2_W_20__5_), .B(_4269__bF_buf4), .Y(_4407_) );
	INVX1 INVX1_134 ( .A(micro_hash_synth_2_W_6__5_), .Y(_4408_) );
	INVX1 INVX1_135 ( .A(micro_hash_synth_2_W_17__5_), .Y(_4409_) );
	OAI21X1 OAI21X1_225 ( .A(_4408_), .B(micro_hash_synth_2_W_11__5_), .C(_4409_), .Y(_4410_) );
	AOI21X1 AOI21X1_100 ( .A(micro_hash_synth_2_W_11__5_), .B(_4408_), .C(_4410_), .Y(_4411_) );
	OAI21X1 OAI21X1_226 ( .A(_4735__bF_buf2), .B(_4411_), .C(_4407_), .Y(_3283_) );
	INVX1 INVX1_136 ( .A(micro_hash_synth_2_W_6__6_), .Y(_4412_) );
	INVX1 INVX1_137 ( .A(micro_hash_synth_2_W_17__6_), .Y(_4413_) );
	OAI21X1 OAI21X1_227 ( .A(_4412_), .B(micro_hash_synth_2_W_11__6_), .C(_4413_), .Y(_4414_) );
	AOI21X1 AOI21X1_101 ( .A(micro_hash_synth_2_W_11__6_), .B(_4412_), .C(_4414_), .Y(_4415_) );
	OAI22X1 OAI22X1_78 ( .A(_4735__bF_buf1), .B(_4415_), .C(_4740__bF_buf2), .D(_4286_), .Y(_3284_) );
	NAND2X1 NAND2X1_158 ( .A(micro_hash_synth_2_W_20__7_), .B(_4269__bF_buf3), .Y(_4416_) );
	INVX1 INVX1_138 ( .A(micro_hash_synth_2_W_17__7_), .Y(_4417_) );
	OAI21X1 OAI21X1_228 ( .A(_4090_), .B(micro_hash_synth_2_W_11__7_), .C(_4417_), .Y(_4418_) );
	AOI21X1 AOI21X1_102 ( .A(micro_hash_synth_2_W_11__7_), .B(_4090_), .C(_4418_), .Y(_4419_) );
	OAI21X1 OAI21X1_229 ( .A(_4735__bF_buf0), .B(_4419_), .C(_4416_), .Y(_3285_) );
	INVX1 INVX1_139 ( .A(bloque_in_1_96_), .Y(_4420_) );
	NAND2X1 NAND2X1_159 ( .A(micro_hash_synth_2_W_12__0_), .B(_4269__bF_buf2), .Y(_4421_) );
	OAI21X1 OAI21X1_230 ( .A(_4420_), .B(_4735__bF_buf15), .C(_4421_), .Y(_3286_) );
	INVX1 INVX1_140 ( .A(bloque_in_1_97_), .Y(_4422_) );
	OAI22X1 OAI22X1_79 ( .A(_4422_), .B(_4735__bF_buf14), .C(_4740__bF_buf1), .D(_4744_), .Y(_3287_) );
	INVX1 INVX1_141 ( .A(bloque_in_1_98_), .Y(_4423_) );
	OAI22X1 OAI22X1_80 ( .A(_4423_), .B(_4735__bF_buf13), .C(_4740__bF_buf0), .D(_4749_), .Y(_3289_) );
	INVX1 INVX1_142 ( .A(bloque_in_1_99_), .Y(_4424_) );
	NAND2X1 NAND2X1_160 ( .A(micro_hash_synth_2_W_12__3_), .B(_4269__bF_buf1), .Y(_4425_) );
	OAI21X1 OAI21X1_231 ( .A(_4424_), .B(_4735__bF_buf12), .C(_4425_), .Y(_3290_) );
	INVX1 INVX1_143 ( .A(bloque_in_1_100_), .Y(_4426_) );
	NAND2X1 NAND2X1_161 ( .A(micro_hash_synth_2_W_12__4_), .B(_4269__bF_buf0), .Y(_4427_) );
	OAI21X1 OAI21X1_232 ( .A(_4426_), .B(_4735__bF_buf11), .C(_4427_), .Y(_3291_) );
	INVX1 INVX1_144 ( .A(bloque_in_1_101_), .Y(_4428_) );
	NAND2X1 NAND2X1_162 ( .A(micro_hash_synth_2_W_12__5_), .B(_4269__bF_buf6), .Y(_4429_) );
	OAI21X1 OAI21X1_233 ( .A(_4428_), .B(_4735__bF_buf10), .C(_4429_), .Y(_3292_) );
	INVX1 INVX1_145 ( .A(bloque_in_1_102_), .Y(_4430_) );
	OAI22X1 OAI22X1_81 ( .A(_4430_), .B(_4735__bF_buf9), .C(_4740__bF_buf13), .D(_4763_), .Y(_3293_) );
	INVX1 INVX1_146 ( .A(bloque_in_1_103_), .Y(_4431_) );
	OAI22X1 OAI22X1_82 ( .A(_4431_), .B(_4735__bF_buf8), .C(_4740__bF_buf12), .D(_4768_), .Y(_3294_) );
	INVX1 INVX1_147 ( .A(micro_hash_synth_2_W_5__0_), .Y(_4432_) );
	OAI21X1 OAI21X1_234 ( .A(_4432_), .B(micro_hash_synth_2_W_10__0_), .C(_3483_), .Y(_4433_) );
	AOI21X1 AOI21X1_103 ( .A(_4432_), .B(micro_hash_synth_2_W_10__0_), .C(_4433_), .Y(_4434_) );
	OAI22X1 OAI22X1_83 ( .A(_4735__bF_buf7), .B(_4434_), .C(_4740__bF_buf11), .D(_4305_), .Y(_3298_) );
	OAI21X1 OAI21X1_235 ( .A(_3555_), .B(micro_hash_synth_2_W_10__1_), .C(_3517_), .Y(_4435_) );
	AOI21X1 AOI21X1_104 ( .A(_3555_), .B(micro_hash_synth_2_W_10__1_), .C(_4435_), .Y(_4436_) );
	OAI22X1 OAI22X1_84 ( .A(_4735__bF_buf6), .B(_4436_), .C(_4740__bF_buf10), .D(_4308_), .Y(_3299_) );
	OAI21X1 OAI21X1_236 ( .A(_3689_), .B(micro_hash_synth_2_W_10__2_), .C(_3618_), .Y(_4437_) );
	AOI21X1 AOI21X1_105 ( .A(_3689_), .B(micro_hash_synth_2_W_10__2_), .C(_4437_), .Y(_4438_) );
	OAI22X1 OAI22X1_85 ( .A(_4735__bF_buf5), .B(_4438_), .C(_4740__bF_buf9), .D(_4311_), .Y(_3300_) );
	INVX1 INVX1_148 ( .A(micro_hash_synth_2_W_5__3_), .Y(_4439_) );
	OAI21X1 OAI21X1_237 ( .A(_4439_), .B(micro_hash_synth_2_W_10__3_), .C(_3748_), .Y(_4440_) );
	AOI21X1 AOI21X1_106 ( .A(_4439_), .B(micro_hash_synth_2_W_10__3_), .C(_4440_), .Y(_4441_) );
	OAI22X1 OAI22X1_86 ( .A(_4735__bF_buf4), .B(_4441_), .C(_4740__bF_buf8), .D(_4315_), .Y(_3301_) );
	INVX1 INVX1_149 ( .A(micro_hash_synth_2_W_5__4_), .Y(_4442_) );
	OAI21X1 OAI21X1_238 ( .A(_4442_), .B(micro_hash_synth_2_W_10__4_), .C(_3845_), .Y(_4443_) );
	AOI21X1 AOI21X1_107 ( .A(_4442_), .B(micro_hash_synth_2_W_10__4_), .C(_4443_), .Y(_4444_) );
	OAI22X1 OAI22X1_87 ( .A(_4735__bF_buf3), .B(_4444_), .C(_4740__bF_buf7), .D(_4319_), .Y(_3303_) );
	INVX1 INVX1_150 ( .A(micro_hash_synth_2_W_5__5_), .Y(_4445_) );
	OAI21X1 OAI21X1_239 ( .A(_4445_), .B(micro_hash_synth_2_W_10__5_), .C(_3902_), .Y(_4446_) );
	AOI21X1 AOI21X1_108 ( .A(_4445_), .B(micro_hash_synth_2_W_10__5_), .C(_4446_), .Y(_4447_) );
	OAI22X1 OAI22X1_88 ( .A(_4735__bF_buf2), .B(_4447_), .C(_4740__bF_buf6), .D(_4323_), .Y(_3304_) );
	INVX1 INVX1_151 ( .A(micro_hash_synth_2_W_5__6_), .Y(_4448_) );
	OAI21X1 OAI21X1_240 ( .A(_4448_), .B(micro_hash_synth_2_W_10__6_), .C(_3985_), .Y(_4449_) );
	AOI21X1 AOI21X1_109 ( .A(_4448_), .B(micro_hash_synth_2_W_10__6_), .C(_4449_), .Y(_4450_) );
	OAI22X1 OAI22X1_89 ( .A(_4735__bF_buf1), .B(_4450_), .C(_4740__bF_buf5), .D(_4327_), .Y(_3305_) );
	INVX1 INVX1_152 ( .A(micro_hash_synth_2_W_5__7_), .Y(_4451_) );
	INVX1 INVX1_153 ( .A(micro_hash_synth_2_W_16__7_), .Y(_4452_) );
	OAI21X1 OAI21X1_241 ( .A(_4451_), .B(micro_hash_synth_2_W_10__7_), .C(_4452_), .Y(_4453_) );
	AOI21X1 AOI21X1_110 ( .A(_4451_), .B(micro_hash_synth_2_W_10__7_), .C(_4453_), .Y(_4454_) );
	OAI22X1 OAI22X1_90 ( .A(_4735__bF_buf0), .B(_4454_), .C(_4740__bF_buf4), .D(_4331_), .Y(_3306_) );
	INVX1 INVX1_154 ( .A(bloque_in_1_40_), .Y(_4455_) );
	OAI22X1 OAI22X1_91 ( .A(_4455_), .B(_4735__bF_buf15), .C(_4740__bF_buf3), .D(_4432_), .Y(_3056_) );
	INVX1 INVX1_155 ( .A(bloque_in_1_41_), .Y(_4456_) );
	OAI22X1 OAI22X1_92 ( .A(_4456_), .B(_4735__bF_buf14), .C(_4740__bF_buf2), .D(_3555_), .Y(_3057_) );
	INVX1 INVX1_156 ( .A(bloque_in_1_42_), .Y(_4457_) );
	OAI22X1 OAI22X1_93 ( .A(_4457_), .B(_4735__bF_buf13), .C(_4740__bF_buf1), .D(_3689_), .Y(_3058_) );
	INVX1 INVX1_157 ( .A(bloque_in_1_43_), .Y(_4458_) );
	OAI22X1 OAI22X1_94 ( .A(_4458_), .B(_4735__bF_buf12), .C(_4740__bF_buf0), .D(_4439_), .Y(_3059_) );
	INVX1 INVX1_158 ( .A(bloque_in_1_44_), .Y(_4459_) );
	OAI22X1 OAI22X1_95 ( .A(_4459_), .B(_4735__bF_buf11), .C(_4740__bF_buf13), .D(_4442_), .Y(_3060_) );
	INVX1 INVX1_159 ( .A(bloque_in_1_45_), .Y(_4460_) );
	OAI22X1 OAI22X1_96 ( .A(_4460_), .B(_4735__bF_buf10), .C(_4740__bF_buf12), .D(_4445_), .Y(_3061_) );
	INVX1 INVX1_160 ( .A(bloque_in_1_46_), .Y(_4461_) );
	OAI22X1 OAI22X1_97 ( .A(_4461_), .B(_4735__bF_buf9), .C(_4740__bF_buf11), .D(_4448_), .Y(_3062_) );
	INVX1 INVX1_161 ( .A(bloque_in_1_47_), .Y(_4462_) );
	OAI22X1 OAI22X1_98 ( .A(_4462_), .B(_4735__bF_buf8), .C(_4740__bF_buf10), .D(_4451_), .Y(_3064_) );
	INVX1 INVX1_162 ( .A(micro_hash_synth_2_W_14__0_), .Y(_4463_) );
	INVX1 INVX1_163 ( .A(bloque_in_1_112_), .Y(_4464_) );
	OAI22X1 OAI22X1_99 ( .A(_4464_), .B(_4735__bF_buf7), .C(_4740__bF_buf9), .D(_4463_), .Y(_3068_) );
	INVX1 INVX1_164 ( .A(micro_hash_synth_2_W_14__1_), .Y(_4465_) );
	INVX1 INVX1_165 ( .A(bloque_in_1_113_), .Y(_4466_) );
	OAI22X1 OAI22X1_100 ( .A(_4466_), .B(_4735__bF_buf6), .C(_4740__bF_buf8), .D(_4465_), .Y(_3069_) );
	INVX1 INVX1_166 ( .A(micro_hash_synth_2_W_14__2_), .Y(_4467_) );
	INVX1 INVX1_167 ( .A(bloque_in_1_114_), .Y(_4468_) );
	OAI22X1 OAI22X1_101 ( .A(_4468_), .B(_4735__bF_buf5), .C(_4740__bF_buf7), .D(_4467_), .Y(_3070_) );
	INVX1 INVX1_168 ( .A(micro_hash_synth_2_W_14__3_), .Y(_4469_) );
	INVX1 INVX1_169 ( .A(bloque_in_1_115_), .Y(_4470_) );
	OAI22X1 OAI22X1_102 ( .A(_4470_), .B(_4735__bF_buf4), .C(_4740__bF_buf6), .D(_4469_), .Y(_3071_) );
	INVX1 INVX1_170 ( .A(micro_hash_synth_2_W_14__4_), .Y(_4471_) );
	INVX1 INVX1_171 ( .A(bloque_in_1_116_), .Y(_4472_) );
	OAI22X1 OAI22X1_103 ( .A(_4472_), .B(_4735__bF_buf3), .C(_4740__bF_buf5), .D(_4471_), .Y(_3072_) );
	INVX1 INVX1_172 ( .A(micro_hash_synth_2_W_14__5_), .Y(_4473_) );
	INVX1 INVX1_173 ( .A(bloque_in_1_117_), .Y(_4474_) );
	OAI22X1 OAI22X1_104 ( .A(_4474_), .B(_4735__bF_buf2), .C(_4740__bF_buf4), .D(_4473_), .Y(_3073_) );
	INVX1 INVX1_174 ( .A(micro_hash_synth_2_W_14__6_), .Y(_4475_) );
	INVX1 INVX1_175 ( .A(bloque_in_1_118_), .Y(_4476_) );
	OAI22X1 OAI22X1_105 ( .A(_4476_), .B(_4735__bF_buf1), .C(_4740__bF_buf3), .D(_4475_), .Y(_3074_) );
	INVX1 INVX1_176 ( .A(micro_hash_synth_2_W_14__7_), .Y(_4477_) );
	INVX1 INVX1_177 ( .A(bloque_in_1_119_), .Y(_4478_) );
	OAI22X1 OAI22X1_106 ( .A(_4478_), .B(_4735__bF_buf0), .C(_4740__bF_buf2), .D(_4477_), .Y(_3075_) );
	INVX1 INVX1_178 ( .A(bloque_in_1_0_), .Y(_4479_) );
	OAI22X1 OAI22X1_107 ( .A(_4479_), .B(_4735__bF_buf15), .C(_4740__bF_buf1), .D(_4841_), .Y(_3077_) );
	INVX1 INVX1_179 ( .A(bloque_in_1_1_), .Y(_4480_) );
	OAI22X1 OAI22X1_108 ( .A(_4480_), .B(_4735__bF_buf14), .C(_4740__bF_buf0), .D(_4842_), .Y(_3078_) );
	INVX1 INVX1_180 ( .A(bloque_in_1_2_), .Y(_4481_) );
	OAI22X1 OAI22X1_109 ( .A(_4481_), .B(_4735__bF_buf13), .C(_4740__bF_buf13), .D(_4843_), .Y(_3080_) );
	INVX1 INVX1_181 ( .A(bloque_in_1_3_), .Y(_4482_) );
	OAI22X1 OAI22X1_110 ( .A(_4482_), .B(_4735__bF_buf12), .C(_4740__bF_buf12), .D(_4844_), .Y(_3081_) );
	INVX1 INVX1_182 ( .A(bloque_in_1_4_), .Y(_4483_) );
	OAI22X1 OAI22X1_111 ( .A(_4483_), .B(_4735__bF_buf11), .C(_4740__bF_buf11), .D(_4845_), .Y(_3082_) );
	INVX1 INVX1_183 ( .A(bloque_in_1_5_), .Y(_4484_) );
	OAI22X1 OAI22X1_112 ( .A(_4484_), .B(_4735__bF_buf10), .C(_4740__bF_buf10), .D(_4846_), .Y(_3083_) );
	INVX1 INVX1_184 ( .A(bloque_in_1_6_), .Y(_4485_) );
	OAI22X1 OAI22X1_113 ( .A(_4485_), .B(_4735__bF_buf9), .C(_4740__bF_buf9), .D(_4847_), .Y(_3084_) );
	INVX1 INVX1_185 ( .A(bloque_in_1_7_), .Y(_4486_) );
	OAI22X1 OAI22X1_114 ( .A(_4486_), .B(_4735__bF_buf8), .C(_4740__bF_buf8), .D(_4848_), .Y(_3085_) );
	INVX1 INVX1_186 ( .A(micro_hash_synth_2_W_15__0_), .Y(_4487_) );
	OAI21X1 OAI21X1_242 ( .A(_4349_), .B(micro_hash_synth_2_W_9__0_), .C(_4487_), .Y(_4488_) );
	AOI21X1 AOI21X1_111 ( .A(_4349_), .B(micro_hash_synth_2_W_9__0_), .C(_4488_), .Y(_4489_) );
	OAI22X1 OAI22X1_115 ( .A(_4735__bF_buf7), .B(_4489_), .C(_4740__bF_buf7), .D(_3480_), .Y(_3086_) );
	INVX1 INVX1_187 ( .A(micro_hash_synth_2_W_15__1_), .Y(_4490_) );
	OAI21X1 OAI21X1_243 ( .A(_4351_), .B(micro_hash_synth_2_W_9__1_), .C(_4490_), .Y(_4491_) );
	AOI21X1 AOI21X1_112 ( .A(_4351_), .B(micro_hash_synth_2_W_9__1_), .C(_4491_), .Y(_4492_) );
	OAI22X1 OAI22X1_116 ( .A(_4735__bF_buf6), .B(_4492_), .C(_4740__bF_buf6), .D(_3513_), .Y(_3087_) );
	INVX1 INVX1_188 ( .A(micro_hash_synth_2_W_15__2_), .Y(_4493_) );
	OAI21X1 OAI21X1_244 ( .A(_4353_), .B(micro_hash_synth_2_W_9__2_), .C(_4493_), .Y(_4494_) );
	AOI21X1 AOI21X1_113 ( .A(_4353_), .B(micro_hash_synth_2_W_9__2_), .C(_4494_), .Y(_4495_) );
	OAI22X1 OAI22X1_117 ( .A(_4735__bF_buf5), .B(_4495_), .C(_4740__bF_buf5), .D(_3614_), .Y(_3088_) );
	INVX1 INVX1_189 ( .A(micro_hash_synth_2_W_15__3_), .Y(_4496_) );
	OAI21X1 OAI21X1_245 ( .A(_4355_), .B(micro_hash_synth_2_W_9__3_), .C(_4496_), .Y(_4497_) );
	AOI21X1 AOI21X1_114 ( .A(_4355_), .B(micro_hash_synth_2_W_9__3_), .C(_4497_), .Y(_4498_) );
	OAI22X1 OAI22X1_118 ( .A(_4735__bF_buf4), .B(_4498_), .C(_4740__bF_buf4), .D(_3744_), .Y(_3089_) );
	INVX1 INVX1_190 ( .A(micro_hash_synth_2_W_15__4_), .Y(_4499_) );
	OAI21X1 OAI21X1_246 ( .A(_4357_), .B(micro_hash_synth_2_W_9__4_), .C(_4499_), .Y(_4500_) );
	AOI21X1 AOI21X1_115 ( .A(_4357_), .B(micro_hash_synth_2_W_9__4_), .C(_4500_), .Y(_4501_) );
	OAI22X1 OAI22X1_119 ( .A(_4735__bF_buf3), .B(_4501_), .C(_4740__bF_buf3), .D(_3841_), .Y(_3090_) );
	INVX1 INVX1_191 ( .A(micro_hash_synth_2_W_15__5_), .Y(_4502_) );
	OAI21X1 OAI21X1_247 ( .A(_4359_), .B(micro_hash_synth_2_W_9__5_), .C(_4502_), .Y(_4503_) );
	AOI21X1 AOI21X1_116 ( .A(_4359_), .B(micro_hash_synth_2_W_9__5_), .C(_4503_), .Y(_4504_) );
	OAI22X1 OAI22X1_120 ( .A(_4735__bF_buf2), .B(_4504_), .C(_4740__bF_buf2), .D(_3898_), .Y(_3091_) );
	OAI21X1 OAI21X1_248 ( .A(_4361_), .B(micro_hash_synth_2_W_9__6_), .C(_4007_), .Y(_4505_) );
	AOI21X1 AOI21X1_117 ( .A(_4361_), .B(micro_hash_synth_2_W_9__6_), .C(_4505_), .Y(_4506_) );
	OAI22X1 OAI22X1_121 ( .A(_4735__bF_buf1), .B(_4506_), .C(_4740__bF_buf1), .D(_3982_), .Y(_3092_) );
	OAI21X1 OAI21X1_249 ( .A(_4363_), .B(micro_hash_synth_2_W_9__7_), .C(_4076_), .Y(_4507_) );
	AOI21X1 AOI21X1_118 ( .A(_4363_), .B(micro_hash_synth_2_W_9__7_), .C(_4507_), .Y(_4508_) );
	OAI22X1 OAI22X1_122 ( .A(_4735__bF_buf0), .B(_4508_), .C(_4740__bF_buf0), .D(_4052_), .Y(_3093_) );
	OAI21X1 OAI21X1_250 ( .A(_4816_), .B(micro_hash_synth_2_W_8__0_), .C(_4463_), .Y(_4509_) );
	AOI21X1 AOI21X1_119 ( .A(micro_hash_synth_2_W_8__0_), .B(_4816_), .C(_4509_), .Y(_4510_) );
	OAI22X1 OAI22X1_123 ( .A(_4735__bF_buf15), .B(_4510_), .C(_4740__bF_buf13), .D(_4384_), .Y(_3094_) );
	OAI21X1 OAI21X1_251 ( .A(_4818_), .B(micro_hash_synth_2_W_8__1_), .C(_4465_), .Y(_4511_) );
	AOI21X1 AOI21X1_120 ( .A(micro_hash_synth_2_W_8__1_), .B(_4818_), .C(_4511_), .Y(_4512_) );
	OAI22X1 OAI22X1_124 ( .A(_4735__bF_buf14), .B(_4512_), .C(_4740__bF_buf12), .D(_4389_), .Y(_3096_) );
	OAI21X1 OAI21X1_252 ( .A(_4820_), .B(micro_hash_synth_2_W_8__2_), .C(_4467_), .Y(_4513_) );
	AOI21X1 AOI21X1_121 ( .A(micro_hash_synth_2_W_8__2_), .B(_4820_), .C(_4513_), .Y(_4514_) );
	OAI22X1 OAI22X1_125 ( .A(_4735__bF_buf13), .B(_4514_), .C(_4740__bF_buf11), .D(_4394_), .Y(_3097_) );
	OAI21X1 OAI21X1_253 ( .A(_4822_), .B(micro_hash_synth_2_W_8__3_), .C(_4469_), .Y(_4515_) );
	AOI21X1 AOI21X1_122 ( .A(micro_hash_synth_2_W_8__3_), .B(_4822_), .C(_4515_), .Y(_4516_) );
	OAI22X1 OAI22X1_126 ( .A(_4735__bF_buf12), .B(_4516_), .C(_4740__bF_buf10), .D(_4399_), .Y(_3098_) );
	OAI21X1 OAI21X1_254 ( .A(_4824_), .B(micro_hash_synth_2_W_8__4_), .C(_4471_), .Y(_4517_) );
	AOI21X1 AOI21X1_123 ( .A(micro_hash_synth_2_W_8__4_), .B(_4824_), .C(_4517_), .Y(_4518_) );
	OAI22X1 OAI22X1_127 ( .A(_4735__bF_buf11), .B(_4518_), .C(_4740__bF_buf9), .D(_4404_), .Y(_3099_) );
	OAI21X1 OAI21X1_255 ( .A(_4826_), .B(micro_hash_synth_2_W_8__5_), .C(_4473_), .Y(_4519_) );
	AOI21X1 AOI21X1_124 ( .A(micro_hash_synth_2_W_8__5_), .B(_4826_), .C(_4519_), .Y(_4520_) );
	OAI22X1 OAI22X1_128 ( .A(_4735__bF_buf10), .B(_4520_), .C(_4740__bF_buf8), .D(_4409_), .Y(_3100_) );
	OAI21X1 OAI21X1_256 ( .A(_4828_), .B(micro_hash_synth_2_W_8__6_), .C(_4475_), .Y(_4521_) );
	AOI21X1 AOI21X1_125 ( .A(micro_hash_synth_2_W_8__6_), .B(_4828_), .C(_4521_), .Y(_4522_) );
	OAI22X1 OAI22X1_129 ( .A(_4735__bF_buf9), .B(_4522_), .C(_4740__bF_buf7), .D(_4413_), .Y(_3101_) );
	OAI21X1 OAI21X1_257 ( .A(_4830_), .B(micro_hash_synth_2_W_8__7_), .C(_4477_), .Y(_4523_) );
	AOI21X1 AOI21X1_126 ( .A(micro_hash_synth_2_W_8__7_), .B(_4830_), .C(_4523_), .Y(_4524_) );
	OAI22X1 OAI22X1_130 ( .A(_4735__bF_buf8), .B(_4524_), .C(_4740__bF_buf6), .D(_4417_), .Y(_3102_) );
	INVX1 INVX1_192 ( .A(bloque_in_1_120_), .Y(_4525_) );
	OAI22X1 OAI22X1_131 ( .A(_4525_), .B(_4735__bF_buf7), .C(_4740__bF_buf5), .D(_4487_), .Y(_3103_) );
	INVX1 INVX1_193 ( .A(bloque_in_1_121_), .Y(_4526_) );
	OAI22X1 OAI22X1_132 ( .A(_4526_), .B(_4735__bF_buf6), .C(_4740__bF_buf4), .D(_4490_), .Y(_3104_) );
	INVX1 INVX1_194 ( .A(bloque_in_1_122_), .Y(_4527_) );
	OAI22X1 OAI22X1_133 ( .A(_4527_), .B(_4735__bF_buf5), .C(_4740__bF_buf3), .D(_4493_), .Y(_3105_) );
	INVX1 INVX1_195 ( .A(bloque_in_1_123_), .Y(_4528_) );
	OAI22X1 OAI22X1_134 ( .A(_4528_), .B(_4735__bF_buf4), .C(_4740__bF_buf2), .D(_4496_), .Y(_3106_) );
	INVX1 INVX1_196 ( .A(bloque_in_1_124_), .Y(_4529_) );
	OAI22X1 OAI22X1_135 ( .A(_4529_), .B(_4735__bF_buf3), .C(_4740__bF_buf1), .D(_4499_), .Y(_3107_) );
	INVX1 INVX1_197 ( .A(bloque_in_1_125_), .Y(_4530_) );
	OAI22X1 OAI22X1_136 ( .A(_4530_), .B(_4735__bF_buf2), .C(_4740__bF_buf0), .D(_4502_), .Y(_3108_) );
	INVX1 INVX1_198 ( .A(bloque_in_1_126_), .Y(_4531_) );
	OAI22X1 OAI22X1_137 ( .A(_4531_), .B(_4735__bF_buf1), .C(_4740__bF_buf13), .D(_4007_), .Y(_3109_) );
	INVX1 INVX1_199 ( .A(bloque_in_1_127_), .Y(_4532_) );
	OAI22X1 OAI22X1_138 ( .A(_4532_), .B(_4735__bF_buf0), .C(_4740__bF_buf12), .D(_4076_), .Y(_3110_) );
	INVX1 INVX1_200 ( .A(bloque_in_1_48_), .Y(_4533_) );
	OAI22X1 OAI22X1_139 ( .A(_4533_), .B(_4735__bF_buf15), .C(_4740__bF_buf11), .D(_4383_), .Y(_3112_) );
	INVX1 INVX1_201 ( .A(bloque_in_1_49_), .Y(_4534_) );
	OAI22X1 OAI22X1_140 ( .A(_4534_), .B(_4735__bF_buf14), .C(_4740__bF_buf10), .D(_4388_), .Y(_3113_) );
	INVX1 INVX1_202 ( .A(bloque_in_1_50_), .Y(_4535_) );
	OAI22X1 OAI22X1_141 ( .A(_4535_), .B(_4735__bF_buf13), .C(_4740__bF_buf9), .D(_4393_), .Y(_3114_) );
	INVX1 INVX1_203 ( .A(bloque_in_1_51_), .Y(_4536_) );
	OAI22X1 OAI22X1_142 ( .A(_4536_), .B(_4735__bF_buf12), .C(_4740__bF_buf8), .D(_4398_), .Y(_3115_) );
	INVX1 INVX1_204 ( .A(bloque_in_1_52_), .Y(_4537_) );
	OAI22X1 OAI22X1_143 ( .A(_4537_), .B(_4735__bF_buf11), .C(_4740__bF_buf7), .D(_4403_), .Y(_3116_) );
	INVX1 INVX1_205 ( .A(bloque_in_1_53_), .Y(_4538_) );
	OAI22X1 OAI22X1_144 ( .A(_4538_), .B(_4735__bF_buf10), .C(_4740__bF_buf6), .D(_4408_), .Y(_3117_) );
	INVX1 INVX1_206 ( .A(bloque_in_1_54_), .Y(_4539_) );
	OAI22X1 OAI22X1_145 ( .A(_4539_), .B(_4735__bF_buf9), .C(_4740__bF_buf5), .D(_4412_), .Y(_3118_) );
	INVX1 INVX1_207 ( .A(bloque_in_1_55_), .Y(_4540_) );
	OAI22X1 OAI22X1_146 ( .A(_4540_), .B(_4735__bF_buf8), .C(_4740__bF_buf4), .D(_4090_), .Y(_3119_) );
	INVX1 INVX1_208 ( .A(micro_hash_synth_2_W_13__0_), .Y(_4541_) );
	INVX1 INVX1_209 ( .A(bloque_in_1_104_), .Y(_4542_) );
	OAI22X1 OAI22X1_147 ( .A(_4542_), .B(_4735__bF_buf7), .C(_4740__bF_buf3), .D(_4541_), .Y(_3120_) );
	INVX1 INVX1_210 ( .A(micro_hash_synth_2_W_13__1_), .Y(_4543_) );
	INVX1 INVX1_211 ( .A(bloque_in_1_105_), .Y(_4544_) );
	OAI22X1 OAI22X1_148 ( .A(_4544_), .B(_4735__bF_buf6), .C(_4740__bF_buf2), .D(_4543_), .Y(_3121_) );
	INVX1 INVX1_212 ( .A(micro_hash_synth_2_W_13__2_), .Y(_4545_) );
	INVX1 INVX1_213 ( .A(bloque_in_1_106_), .Y(_4546_) );
	OAI22X1 OAI22X1_149 ( .A(_4546_), .B(_4735__bF_buf5), .C(_4740__bF_buf1), .D(_4545_), .Y(_3122_) );
	INVX1 INVX1_214 ( .A(micro_hash_synth_2_W_13__3_), .Y(_4547_) );
	INVX1 INVX1_215 ( .A(bloque_in_1_107_), .Y(_4548_) );
	OAI22X1 OAI22X1_150 ( .A(_4548_), .B(_4735__bF_buf4), .C(_4740__bF_buf0), .D(_4547_), .Y(_3123_) );
	INVX1 INVX1_216 ( .A(micro_hash_synth_2_W_13__4_), .Y(_4549_) );
	INVX1 INVX1_217 ( .A(bloque_in_1_108_), .Y(_4550_) );
	OAI22X1 OAI22X1_151 ( .A(_4550_), .B(_4735__bF_buf3), .C(_4740__bF_buf13), .D(_4549_), .Y(_3124_) );
	INVX1 INVX1_218 ( .A(micro_hash_synth_2_W_13__5_), .Y(_4551_) );
	INVX1 INVX1_219 ( .A(bloque_in_1_109_), .Y(_4552_) );
	OAI22X1 OAI22X1_152 ( .A(_4552_), .B(_4735__bF_buf2), .C(_4740__bF_buf12), .D(_4551_), .Y(_3125_) );
	INVX1 INVX1_220 ( .A(micro_hash_synth_2_W_13__6_), .Y(_4553_) );
	INVX1 INVX1_221 ( .A(bloque_in_1_110_), .Y(_4554_) );
	OAI22X1 OAI22X1_153 ( .A(_4554_), .B(_4735__bF_buf1), .C(_4740__bF_buf11), .D(_4553_), .Y(_3126_) );
	INVX1 INVX1_222 ( .A(micro_hash_synth_2_W_13__7_), .Y(_4555_) );
	INVX1 INVX1_223 ( .A(bloque_in_1_111_), .Y(_4556_) );
	OAI22X1 OAI22X1_154 ( .A(_4556_), .B(_4735__bF_buf0), .C(_4740__bF_buf10), .D(_4555_), .Y(_3128_) );
	OAI21X1 OAI21X1_258 ( .A(_4849_), .B(micro_hash_synth_2_W_7__0_), .C(_4541_), .Y(_4557_) );
	AOI21X1 AOI21X1_127 ( .A(_4849_), .B(micro_hash_synth_2_W_7__0_), .C(_4557_), .Y(_4558_) );
	OAI22X1 OAI22X1_155 ( .A(_4735__bF_buf15), .B(_4558_), .C(_4740__bF_buf9), .D(_3483_), .Y(_3129_) );
	OAI21X1 OAI21X1_259 ( .A(_4850_), .B(micro_hash_synth_2_W_7__1_), .C(_4543_), .Y(_4559_) );
	AOI21X1 AOI21X1_128 ( .A(_4850_), .B(micro_hash_synth_2_W_7__1_), .C(_4559_), .Y(_4560_) );
	OAI22X1 OAI22X1_156 ( .A(_4735__bF_buf14), .B(_4560_), .C(_4740__bF_buf8), .D(_3517_), .Y(_3130_) );
	OAI21X1 OAI21X1_260 ( .A(_4851_), .B(micro_hash_synth_2_W_7__2_), .C(_4545_), .Y(_4561_) );
	AOI21X1 AOI21X1_129 ( .A(_4851_), .B(micro_hash_synth_2_W_7__2_), .C(_4561_), .Y(_4562_) );
	OAI22X1 OAI22X1_157 ( .A(_4735__bF_buf13), .B(_4562_), .C(_4740__bF_buf7), .D(_3618_), .Y(_3131_) );
	OAI21X1 OAI21X1_261 ( .A(_4852_), .B(micro_hash_synth_2_W_7__3_), .C(_4547_), .Y(_4563_) );
	AOI21X1 AOI21X1_130 ( .A(_4852_), .B(micro_hash_synth_2_W_7__3_), .C(_4563_), .Y(_4564_) );
	OAI22X1 OAI22X1_158 ( .A(_4735__bF_buf12), .B(_4564_), .C(_4740__bF_buf6), .D(_3748_), .Y(_3132_) );
	OAI21X1 OAI21X1_262 ( .A(_4853_), .B(micro_hash_synth_2_W_7__4_), .C(_4549_), .Y(_4565_) );
	AOI21X1 AOI21X1_131 ( .A(_4853_), .B(micro_hash_synth_2_W_7__4_), .C(_4565_), .Y(_4566_) );
	OAI22X1 OAI22X1_159 ( .A(_4735__bF_buf11), .B(_4566_), .C(_4740__bF_buf5), .D(_3845_), .Y(_3133_) );
	OAI21X1 OAI21X1_263 ( .A(_4854_), .B(micro_hash_synth_2_W_7__5_), .C(_4551_), .Y(_4567_) );
	AOI21X1 AOI21X1_132 ( .A(_4854_), .B(micro_hash_synth_2_W_7__5_), .C(_4567_), .Y(_4568_) );
	OAI22X1 OAI22X1_160 ( .A(_4735__bF_buf10), .B(_4568_), .C(_4740__bF_buf4), .D(_3902_), .Y(_3134_) );
	OAI21X1 OAI21X1_264 ( .A(_4855_), .B(micro_hash_synth_2_W_7__6_), .C(_4553_), .Y(_4569_) );
	AOI21X1 AOI21X1_133 ( .A(_4855_), .B(micro_hash_synth_2_W_7__6_), .C(_4569_), .Y(_4570_) );
	OAI22X1 OAI22X1_161 ( .A(_4735__bF_buf9), .B(_4570_), .C(_4740__bF_buf3), .D(_3985_), .Y(_3135_) );
	OAI21X1 OAI21X1_265 ( .A(_4856_), .B(micro_hash_synth_2_W_7__7_), .C(_4555_), .Y(_4571_) );
	AOI21X1 AOI21X1_134 ( .A(_4856_), .B(micro_hash_synth_2_W_7__7_), .C(_4571_), .Y(_4572_) );
	OAI22X1 OAI22X1_162 ( .A(_4735__bF_buf8), .B(_4572_), .C(_4740__bF_buf2), .D(_4452_), .Y(_3136_) );
	INVX1 INVX1_224 ( .A(bloque_in_1_8_), .Y(_4573_) );
	OAI22X1 OAI22X1_163 ( .A(_4573_), .B(_4735__bF_buf7), .C(_4740__bF_buf1), .D(_4833_), .Y(_3137_) );
	INVX1 INVX1_225 ( .A(bloque_in_1_9_), .Y(_4574_) );
	OAI22X1 OAI22X1_164 ( .A(_4574_), .B(_4735__bF_buf6), .C(_4740__bF_buf0), .D(_4834_), .Y(_3138_) );
	INVX1 INVX1_226 ( .A(bloque_in_1_10_), .Y(_4575_) );
	OAI22X1 OAI22X1_165 ( .A(_4575_), .B(_4735__bF_buf5), .C(_4740__bF_buf13), .D(_4835_), .Y(_3139_) );
	INVX1 INVX1_227 ( .A(bloque_in_1_11_), .Y(_4576_) );
	OAI22X1 OAI22X1_166 ( .A(_4576_), .B(_4735__bF_buf4), .C(_4740__bF_buf12), .D(_4836_), .Y(_3140_) );
	INVX1 INVX1_228 ( .A(bloque_in_1_12_), .Y(_4577_) );
	OAI22X1 OAI22X1_167 ( .A(_4577_), .B(_4735__bF_buf3), .C(_4740__bF_buf11), .D(_4837_), .Y(_3141_) );
	INVX1 INVX1_229 ( .A(bloque_in_1_13_), .Y(_4578_) );
	OAI22X1 OAI22X1_168 ( .A(_4578_), .B(_4735__bF_buf2), .C(_4740__bF_buf10), .D(_4838_), .Y(_3142_) );
	INVX1 INVX1_230 ( .A(bloque_in_1_14_), .Y(_4579_) );
	OAI22X1 OAI22X1_169 ( .A(_4579_), .B(_4735__bF_buf1), .C(_4740__bF_buf9), .D(_4839_), .Y(_3144_) );
	INVX1 INVX1_231 ( .A(bloque_in_1_15_), .Y(_4580_) );
	OAI22X1 OAI22X1_170 ( .A(_4580_), .B(_4735__bF_buf0), .C(_4740__bF_buf8), .D(_4840_), .Y(_3145_) );
	INVX1 INVX1_232 ( .A(bloque_in_1_80_), .Y(_4581_) );
	NAND2X1 NAND2X1_163 ( .A(micro_hash_synth_2_W_10__0_), .B(_4269__bF_buf5), .Y(_4582_) );
	OAI21X1 OAI21X1_266 ( .A(_4581_), .B(_4735__bF_buf15), .C(_4582_), .Y(_3146_) );
	INVX1 INVX1_233 ( .A(bloque_in_1_81_), .Y(_4583_) );
	OAI22X1 OAI22X1_171 ( .A(_4583_), .B(_4735__bF_buf14), .C(_4740__bF_buf7), .D(_3546_), .Y(_3147_) );
	INVX1 INVX1_234 ( .A(bloque_in_1_82_), .Y(_4584_) );
	OAI22X1 OAI22X1_172 ( .A(_4584_), .B(_4735__bF_buf13), .C(_4740__bF_buf6), .D(_3646_), .Y(_3148_) );
	INVX1 INVX1_235 ( .A(bloque_in_1_83_), .Y(_4585_) );
	OAI22X1 OAI22X1_173 ( .A(_4585_), .B(_4735__bF_buf12), .C(_4740__bF_buf5), .D(_3761_), .Y(_3149_) );
	INVX1 INVX1_236 ( .A(bloque_in_1_84_), .Y(_4586_) );
	OAI22X1 OAI22X1_174 ( .A(_4586_), .B(_4735__bF_buf11), .C(_4740__bF_buf4), .D(_3827_), .Y(_3150_) );
	INVX1 INVX1_237 ( .A(bloque_in_1_85_), .Y(_4587_) );
	OAI22X1 OAI22X1_175 ( .A(_4587_), .B(_4735__bF_buf10), .C(_4740__bF_buf3), .D(_3929_), .Y(_3151_) );
	INVX1 INVX1_238 ( .A(bloque_in_1_86_), .Y(_4588_) );
	OAI22X1 OAI22X1_176 ( .A(_4588_), .B(_4735__bF_buf9), .C(_4740__bF_buf2), .D(_4015_), .Y(_3152_) );
	INVX1 INVX1_239 ( .A(bloque_in_1_87_), .Y(_4589_) );
	OAI22X1 OAI22X1_177 ( .A(_4589_), .B(_4735__bF_buf8), .C(_4740__bF_buf1), .D(_4265_), .Y(_3153_) );
	INVX1 INVX1_240 ( .A(bloque_in_1_88_), .Y(_4590_) );
	NAND2X1 NAND2X1_164 ( .A(micro_hash_synth_2_W_11__0_), .B(_4269__bF_buf4), .Y(_4591_) );
	OAI21X1 OAI21X1_267 ( .A(_4590_), .B(_4735__bF_buf7), .C(_4591_), .Y(_3154_) );
	INVX1 INVX1_241 ( .A(bloque_in_1_89_), .Y(_4592_) );
	OAI22X1 OAI22X1_178 ( .A(_4592_), .B(_4735__bF_buf6), .C(_4740__bF_buf0), .D(_4776_), .Y(_3155_) );
	INVX1 INVX1_242 ( .A(bloque_in_1_90_), .Y(_4593_) );
	OAI22X1 OAI22X1_179 ( .A(_4593_), .B(_4735__bF_buf5), .C(_4740__bF_buf13), .D(_4781_), .Y(_3156_) );
	INVX1 INVX1_243 ( .A(bloque_in_1_91_), .Y(_4594_) );
	NAND2X1 NAND2X1_165 ( .A(micro_hash_synth_2_W_11__3_), .B(_4269__bF_buf3), .Y(_4595_) );
	OAI21X1 OAI21X1_268 ( .A(_4594_), .B(_4735__bF_buf4), .C(_4595_), .Y(_3157_) );
	INVX1 INVX1_244 ( .A(bloque_in_1_92_), .Y(_4596_) );
	NAND2X1 NAND2X1_166 ( .A(micro_hash_synth_2_W_11__4_), .B(_4269__bF_buf2), .Y(_4597_) );
	OAI21X1 OAI21X1_269 ( .A(_4596_), .B(_4735__bF_buf3), .C(_4597_), .Y(_3158_) );
	INVX1 INVX1_245 ( .A(bloque_in_1_93_), .Y(_4598_) );
	NAND2X1 NAND2X1_167 ( .A(micro_hash_synth_2_W_11__5_), .B(_4269__bF_buf1), .Y(_4599_) );
	OAI21X1 OAI21X1_270 ( .A(_4598_), .B(_4735__bF_buf2), .C(_4599_), .Y(_3159_) );
	INVX1 INVX1_246 ( .A(bloque_in_1_94_), .Y(_4600_) );
	NAND2X1 NAND2X1_168 ( .A(micro_hash_synth_2_W_11__6_), .B(_4269__bF_buf0), .Y(_4601_) );
	OAI21X1 OAI21X1_271 ( .A(_4600_), .B(_4735__bF_buf1), .C(_4601_), .Y(_3160_) );
	INVX1 INVX1_247 ( .A(bloque_in_1_95_), .Y(_4602_) );
	NAND2X1 NAND2X1_169 ( .A(micro_hash_synth_2_W_11__7_), .B(_4269__bF_buf6), .Y(_4603_) );
	OAI21X1 OAI21X1_272 ( .A(_4602_), .B(_4735__bF_buf0), .C(_4603_), .Y(_3161_) );
	INVX1 INVX1_248 ( .A(bloque_in_1_16_), .Y(_4604_) );
	OAI22X1 OAI22X1_180 ( .A(_4604_), .B(_4735__bF_buf15), .C(_4740__bF_buf12), .D(_4849_), .Y(_3162_) );
	INVX1 INVX1_249 ( .A(bloque_in_1_17_), .Y(_4605_) );
	OAI22X1 OAI22X1_181 ( .A(_4605_), .B(_4735__bF_buf14), .C(_4740__bF_buf11), .D(_4850_), .Y(_3163_) );
	INVX1 INVX1_250 ( .A(bloque_in_1_18_), .Y(_4606_) );
	OAI22X1 OAI22X1_182 ( .A(_4606_), .B(_4735__bF_buf13), .C(_4740__bF_buf10), .D(_4851_), .Y(_3164_) );
	INVX1 INVX1_251 ( .A(bloque_in_1_19_), .Y(_4607_) );
	OAI22X1 OAI22X1_183 ( .A(_4607_), .B(_4735__bF_buf12), .C(_4740__bF_buf9), .D(_4852_), .Y(_3165_) );
	INVX1 INVX1_252 ( .A(bloque_in_1_20_), .Y(_4608_) );
	OAI22X1 OAI22X1_184 ( .A(_4608_), .B(_4735__bF_buf11), .C(_4740__bF_buf8), .D(_4853_), .Y(_3166_) );
	INVX1 INVX1_253 ( .A(bloque_in_1_21_), .Y(_4609_) );
	OAI22X1 OAI22X1_185 ( .A(_4609_), .B(_4735__bF_buf10), .C(_4740__bF_buf7), .D(_4854_), .Y(_3167_) );
	INVX1 INVX1_254 ( .A(bloque_in_1_22_), .Y(_4610_) );
	OAI22X1 OAI22X1_186 ( .A(_4610_), .B(_4735__bF_buf9), .C(_4740__bF_buf6), .D(_4855_), .Y(_3168_) );
	INVX1 INVX1_255 ( .A(bloque_in_1_23_), .Y(_4611_) );
	OAI22X1 OAI22X1_187 ( .A(_4611_), .B(_4735__bF_buf8), .C(_4740__bF_buf5), .D(_4856_), .Y(_3169_) );
	INVX1 INVX1_256 ( .A(micro_hash_synth_2_W_27__0_), .Y(_4612_) );
	OAI21X1 OAI21X1_273 ( .A(_4541_), .B(micro_hash_synth_2_W_18__0_), .C(_4244_), .Y(_4613_) );
	AOI21X1 AOI21X1_135 ( .A(_4541_), .B(micro_hash_synth_2_W_18__0_), .C(_4613_), .Y(_4614_) );
	OAI22X1 OAI22X1_188 ( .A(_4735__bF_buf7), .B(_4614_), .C(_4740__bF_buf4), .D(_4612_), .Y(_3170_) );
	INVX1 INVX1_257 ( .A(micro_hash_synth_2_W_27__1_), .Y(_4615_) );
	OAI21X1 OAI21X1_274 ( .A(_4543_), .B(micro_hash_synth_2_W_18__1_), .C(_3533_), .Y(_4616_) );
	AOI21X1 AOI21X1_136 ( .A(_4543_), .B(micro_hash_synth_2_W_18__1_), .C(_4616_), .Y(_4617_) );
	OAI22X1 OAI22X1_189 ( .A(_4735__bF_buf6), .B(_4617_), .C(_4740__bF_buf3), .D(_4615_), .Y(_3171_) );
	INVX1 INVX1_258 ( .A(micro_hash_synth_2_W_27__2_), .Y(_4618_) );
	OAI21X1 OAI21X1_275 ( .A(_4545_), .B(micro_hash_synth_2_W_18__2_), .C(_3629_), .Y(_4619_) );
	AOI21X1 AOI21X1_137 ( .A(_4545_), .B(micro_hash_synth_2_W_18__2_), .C(_4619_), .Y(_4620_) );
	OAI22X1 OAI22X1_190 ( .A(_4735__bF_buf5), .B(_4620_), .C(_4740__bF_buf2), .D(_4618_), .Y(_3172_) );
	INVX1 INVX1_259 ( .A(micro_hash_synth_2_W_27__3_), .Y(_4621_) );
	OAI21X1 OAI21X1_276 ( .A(_4547_), .B(micro_hash_synth_2_W_18__3_), .C(_3729_), .Y(_4622_) );
	AOI21X1 AOI21X1_138 ( .A(_4547_), .B(micro_hash_synth_2_W_18__3_), .C(_4622_), .Y(_4623_) );
	OAI22X1 OAI22X1_191 ( .A(_4735__bF_buf4), .B(_4623_), .C(_4740__bF_buf1), .D(_4621_), .Y(_3173_) );
	INVX1 INVX1_260 ( .A(micro_hash_synth_2_W_27__4_), .Y(_4624_) );
	OAI21X1 OAI21X1_277 ( .A(_4549_), .B(micro_hash_synth_2_W_18__4_), .C(_3813_), .Y(_4625_) );
	AOI21X1 AOI21X1_139 ( .A(_4549_), .B(micro_hash_synth_2_W_18__4_), .C(_4625_), .Y(_4626_) );
	OAI22X1 OAI22X1_192 ( .A(_4735__bF_buf3), .B(_4626_), .C(_4740__bF_buf0), .D(_4624_), .Y(_3174_) );
	INVX1 INVX1_261 ( .A(micro_hash_synth_2_W_27__5_), .Y(_4627_) );
	OAI21X1 OAI21X1_278 ( .A(_4551_), .B(micro_hash_synth_2_W_18__5_), .C(_3915_), .Y(_4628_) );
	AOI21X1 AOI21X1_140 ( .A(_4551_), .B(micro_hash_synth_2_W_18__5_), .C(_4628_), .Y(_4629_) );
	OAI22X1 OAI22X1_193 ( .A(_4735__bF_buf2), .B(_4629_), .C(_4740__bF_buf13), .D(_4627_), .Y(_3175_) );
	INVX1 INVX1_262 ( .A(micro_hash_synth_2_W_27__6_), .Y(_4630_) );
	OAI21X1 OAI21X1_279 ( .A(_4553_), .B(micro_hash_synth_2_W_18__6_), .C(_3996_), .Y(_4631_) );
	AOI21X1 AOI21X1_141 ( .A(_4553_), .B(micro_hash_synth_2_W_18__6_), .C(_4631_), .Y(_4632_) );
	OAI22X1 OAI22X1_194 ( .A(_4735__bF_buf1), .B(_4632_), .C(_4740__bF_buf12), .D(_4630_), .Y(_3176_) );
	INVX1 INVX1_263 ( .A(micro_hash_synth_2_W_27__7_), .Y(_4633_) );
	OAI21X1 OAI21X1_280 ( .A(_4555_), .B(micro_hash_synth_2_W_18__7_), .C(_4068_), .Y(_4634_) );
	AOI21X1 AOI21X1_142 ( .A(_4555_), .B(micro_hash_synth_2_W_18__7_), .C(_4634_), .Y(_4635_) );
	OAI22X1 OAI22X1_195 ( .A(_4735__bF_buf0), .B(_4635_), .C(_4740__bF_buf11), .D(_4633_), .Y(_3177_) );
	INVX1 INVX1_264 ( .A(micro_hash_synth_2_W_28__0_), .Y(_4636_) );
	OAI21X1 OAI21X1_281 ( .A(_4463_), .B(micro_hash_synth_2_W_19__0_), .C(_4772_), .Y(_4637_) );
	AOI21X1 AOI21X1_143 ( .A(_4463_), .B(micro_hash_synth_2_W_19__0_), .C(_4637_), .Y(_4638_) );
	OAI22X1 OAI22X1_196 ( .A(_4735__bF_buf15), .B(_4638_), .C(_4740__bF_buf10), .D(_4636_), .Y(_3178_) );
	INVX1 INVX1_265 ( .A(micro_hash_synth_2_W_28__1_), .Y(_4639_) );
	OAI21X1 OAI21X1_282 ( .A(_4465_), .B(micro_hash_synth_2_W_19__1_), .C(_4775_), .Y(_4640_) );
	AOI21X1 AOI21X1_144 ( .A(_4465_), .B(micro_hash_synth_2_W_19__1_), .C(_4640_), .Y(_4641_) );
	OAI22X1 OAI22X1_197 ( .A(_4735__bF_buf14), .B(_4641_), .C(_4740__bF_buf9), .D(_4639_), .Y(_3179_) );
	INVX1 INVX1_266 ( .A(micro_hash_synth_2_W_28__2_), .Y(_4642_) );
	OAI21X1 OAI21X1_283 ( .A(_4467_), .B(micro_hash_synth_2_W_19__2_), .C(_4780_), .Y(_4643_) );
	AOI21X1 AOI21X1_145 ( .A(_4467_), .B(micro_hash_synth_2_W_19__2_), .C(_4643_), .Y(_4644_) );
	OAI22X1 OAI22X1_198 ( .A(_4735__bF_buf13), .B(_4644_), .C(_4740__bF_buf8), .D(_4642_), .Y(_3180_) );
	INVX1 INVX1_267 ( .A(micro_hash_synth_2_W_28__3_), .Y(_4645_) );
	OAI21X1 OAI21X1_284 ( .A(_4469_), .B(micro_hash_synth_2_W_19__3_), .C(_4785_), .Y(_4646_) );
	AOI21X1 AOI21X1_146 ( .A(_4469_), .B(micro_hash_synth_2_W_19__3_), .C(_4646_), .Y(_4647_) );
	OAI22X1 OAI22X1_199 ( .A(_4735__bF_buf12), .B(_4647_), .C(_4740__bF_buf7), .D(_4645_), .Y(_3181_) );
	INVX1 INVX1_268 ( .A(micro_hash_synth_2_W_28__4_), .Y(_4648_) );
	OAI21X1 OAI21X1_285 ( .A(_4471_), .B(micro_hash_synth_2_W_19__4_), .C(_4788_), .Y(_4649_) );
	AOI21X1 AOI21X1_147 ( .A(_4471_), .B(micro_hash_synth_2_W_19__4_), .C(_4649_), .Y(_4650_) );
	OAI22X1 OAI22X1_200 ( .A(_4735__bF_buf11), .B(_4650_), .C(_4740__bF_buf6), .D(_4648_), .Y(_3182_) );
	INVX1 INVX1_269 ( .A(micro_hash_synth_2_W_28__5_), .Y(_4651_) );
	OAI21X1 OAI21X1_286 ( .A(_4473_), .B(micro_hash_synth_2_W_19__5_), .C(_4791_), .Y(_4652_) );
	AOI21X1 AOI21X1_148 ( .A(_4473_), .B(micro_hash_synth_2_W_19__5_), .C(_4652_), .Y(_4653_) );
	OAI22X1 OAI22X1_201 ( .A(_4735__bF_buf10), .B(_4653_), .C(_4740__bF_buf5), .D(_4651_), .Y(_3183_) );
	INVX1 INVX1_270 ( .A(micro_hash_synth_2_W_28__6_), .Y(_4654_) );
	OAI21X1 OAI21X1_287 ( .A(_4475_), .B(micro_hash_synth_2_W_19__6_), .C(_4794_), .Y(_4655_) );
	AOI21X1 AOI21X1_149 ( .A(_4475_), .B(micro_hash_synth_2_W_19__6_), .C(_4655_), .Y(_4656_) );
	OAI22X1 OAI22X1_202 ( .A(_4735__bF_buf9), .B(_4656_), .C(_4740__bF_buf4), .D(_4654_), .Y(_3184_) );
	INVX1 INVX1_271 ( .A(micro_hash_synth_2_W_28__7_), .Y(_4657_) );
	OAI21X1 OAI21X1_288 ( .A(_4477_), .B(micro_hash_synth_2_W_19__7_), .C(_4797_), .Y(_4658_) );
	AOI21X1 AOI21X1_150 ( .A(_4477_), .B(micro_hash_synth_2_W_19__7_), .C(_4658_), .Y(_4659_) );
	OAI22X1 OAI22X1_203 ( .A(_4735__bF_buf8), .B(_4659_), .C(_4740__bF_buf3), .D(_4657_), .Y(_3185_) );
	NAND2X1 NAND2X1_170 ( .A(micro_hash_synth_2_W_29__0_), .B(_4269__bF_buf5), .Y(_4660_) );
	OAI21X1 OAI21X1_289 ( .A(_4487_), .B(micro_hash_synth_2_W_20__0_), .C(_4728_), .Y(_4661_) );
	AOI21X1 AOI21X1_151 ( .A(_4487_), .B(micro_hash_synth_2_W_20__0_), .C(_4661_), .Y(_4662_) );
	OAI21X1 OAI21X1_290 ( .A(_4735__bF_buf7), .B(_4662_), .C(_4660_), .Y(_3186_) );
	OAI21X1 OAI21X1_291 ( .A(_4490_), .B(micro_hash_synth_2_W_20__1_), .C(_4743_), .Y(_4663_) );
	AOI21X1 AOI21X1_152 ( .A(_4490_), .B(micro_hash_synth_2_W_20__1_), .C(_4663_), .Y(_4664_) );
	OAI22X1 OAI22X1_204 ( .A(_4735__bF_buf6), .B(_4664_), .C(_4740__bF_buf2), .D(_3524_), .Y(_3187_) );
	OAI21X1 OAI21X1_292 ( .A(_4493_), .B(micro_hash_synth_2_W_20__2_), .C(_4748_), .Y(_4665_) );
	AOI21X1 AOI21X1_153 ( .A(_4493_), .B(micro_hash_synth_2_W_20__2_), .C(_4665_), .Y(_4666_) );
	OAI22X1 OAI22X1_205 ( .A(_4735__bF_buf5), .B(_4666_), .C(_4740__bF_buf1), .D(_3674_), .Y(_3188_) );
	NAND2X1 NAND2X1_171 ( .A(micro_hash_synth_2_W_29__3_), .B(_4269__bF_buf4), .Y(_4667_) );
	OAI21X1 OAI21X1_293 ( .A(_4496_), .B(micro_hash_synth_2_W_20__3_), .C(_4753_), .Y(_4668_) );
	AOI21X1 AOI21X1_154 ( .A(_4496_), .B(micro_hash_synth_2_W_20__3_), .C(_4668_), .Y(_4669_) );
	OAI21X1 OAI21X1_294 ( .A(_4735__bF_buf4), .B(_4669_), .C(_4667_), .Y(_3189_) );
	NAND2X1 NAND2X1_172 ( .A(micro_hash_synth_2_W_29__4_), .B(_4269__bF_buf3), .Y(_4670_) );
	OAI21X1 OAI21X1_295 ( .A(_4499_), .B(micro_hash_synth_2_W_20__4_), .C(_4756_), .Y(_4671_) );
	AOI21X1 AOI21X1_155 ( .A(_4499_), .B(micro_hash_synth_2_W_20__4_), .C(_4671_), .Y(_4672_) );
	OAI21X1 OAI21X1_296 ( .A(_4735__bF_buf3), .B(_4672_), .C(_4670_), .Y(_3190_) );
	NAND2X1 NAND2X1_173 ( .A(micro_hash_synth_2_W_29__5_), .B(_4269__bF_buf2), .Y(_4673_) );
	OAI21X1 OAI21X1_297 ( .A(_4502_), .B(micro_hash_synth_2_W_20__5_), .C(_4759_), .Y(_4674_) );
	AOI21X1 AOI21X1_156 ( .A(_4502_), .B(micro_hash_synth_2_W_20__5_), .C(_4674_), .Y(_4675_) );
	OAI21X1 OAI21X1_298 ( .A(_4735__bF_buf2), .B(_4675_), .C(_4673_), .Y(_3191_) );
	NAND2X1 NAND2X1_174 ( .A(micro_hash_synth_2_W_29__6_), .B(_4269__bF_buf1), .Y(_4676_) );
	OAI21X1 OAI21X1_299 ( .A(_4007_), .B(micro_hash_synth_2_W_20__6_), .C(_4762_), .Y(_4677_) );
	AOI21X1 AOI21X1_157 ( .A(_4007_), .B(micro_hash_synth_2_W_20__6_), .C(_4677_), .Y(_4678_) );
	OAI21X1 OAI21X1_300 ( .A(_4735__bF_buf1), .B(_4678_), .C(_4676_), .Y(_3192_) );
	NAND2X1 NAND2X1_175 ( .A(micro_hash_synth_2_W_29__7_), .B(_4269__bF_buf0), .Y(_4679_) );
	OAI21X1 OAI21X1_301 ( .A(_4076_), .B(micro_hash_synth_2_W_20__7_), .C(_4767_), .Y(_4680_) );
	AOI21X1 AOI21X1_158 ( .A(_4076_), .B(micro_hash_synth_2_W_20__7_), .C(_4680_), .Y(_4681_) );
	OAI21X1 OAI21X1_302 ( .A(_4735__bF_buf0), .B(_4681_), .C(_4679_), .Y(_3193_) );
	NAND2X1 NAND2X1_176 ( .A(micro_hash_synth_2_W_30__0_), .B(_4269__bF_buf6), .Y(_4682_) );
	OAI21X1 OAI21X1_303 ( .A(_3483_), .B(micro_hash_synth_2_W_21__0_), .C(_4612_), .Y(_4683_) );
	AOI21X1 AOI21X1_159 ( .A(_3483_), .B(micro_hash_synth_2_W_21__0_), .C(_4683_), .Y(_4684_) );
	OAI21X1 OAI21X1_304 ( .A(_4735__bF_buf15), .B(_4684_), .C(_4682_), .Y(_3194_) );
	NAND2X1 NAND2X1_177 ( .A(micro_hash_synth_2_W_30__1_), .B(_4269__bF_buf5), .Y(_4685_) );
	OAI21X1 OAI21X1_305 ( .A(_3517_), .B(micro_hash_synth_2_W_21__1_), .C(_4615_), .Y(_4686_) );
	AOI21X1 AOI21X1_160 ( .A(_3517_), .B(micro_hash_synth_2_W_21__1_), .C(_4686_), .Y(_4687_) );
	OAI21X1 OAI21X1_306 ( .A(_4735__bF_buf14), .B(_4687_), .C(_4685_), .Y(_3195_) );
	NAND2X1 NAND2X1_178 ( .A(micro_hash_synth_2_W_30__2_), .B(_4269__bF_buf4), .Y(_4688_) );
	OAI21X1 OAI21X1_307 ( .A(_3618_), .B(micro_hash_synth_2_W_21__2_), .C(_4618_), .Y(_4689_) );
	AOI21X1 AOI21X1_161 ( .A(_3618_), .B(micro_hash_synth_2_W_21__2_), .C(_4689_), .Y(_4690_) );
	OAI21X1 OAI21X1_308 ( .A(_4735__bF_buf13), .B(_4690_), .C(_4688_), .Y(_3196_) );
	NAND2X1 NAND2X1_179 ( .A(micro_hash_synth_2_W_30__3_), .B(_4269__bF_buf3), .Y(_4691_) );
	OAI21X1 OAI21X1_309 ( .A(_3748_), .B(micro_hash_synth_2_W_21__3_), .C(_4621_), .Y(_4692_) );
	AOI21X1 AOI21X1_162 ( .A(_3748_), .B(micro_hash_synth_2_W_21__3_), .C(_4692_), .Y(_4693_) );
	OAI21X1 OAI21X1_310 ( .A(_4735__bF_buf12), .B(_4693_), .C(_4691_), .Y(_3197_) );
	NAND2X1 NAND2X1_180 ( .A(micro_hash_synth_2_W_30__4_), .B(_4269__bF_buf2), .Y(_4694_) );
	OAI21X1 OAI21X1_311 ( .A(_3845_), .B(micro_hash_synth_2_W_21__4_), .C(_4624_), .Y(_4695_) );
	AOI21X1 AOI21X1_163 ( .A(_3845_), .B(micro_hash_synth_2_W_21__4_), .C(_4695_), .Y(_4696_) );
	OAI21X1 OAI21X1_312 ( .A(_4735__bF_buf11), .B(_4696_), .C(_4694_), .Y(_3198_) );
	NAND2X1 NAND2X1_181 ( .A(micro_hash_synth_2_W_30__5_), .B(_4269__bF_buf1), .Y(_4697_) );
	OAI21X1 OAI21X1_313 ( .A(_3902_), .B(micro_hash_synth_2_W_21__5_), .C(_4627_), .Y(_4698_) );
	AOI21X1 AOI21X1_164 ( .A(_3902_), .B(micro_hash_synth_2_W_21__5_), .C(_4698_), .Y(_4699_) );
	OAI21X1 OAI21X1_314 ( .A(_4735__bF_buf10), .B(_4699_), .C(_4697_), .Y(_3199_) );
	NAND2X1 NAND2X1_182 ( .A(micro_hash_synth_2_W_30__6_), .B(_4269__bF_buf0), .Y(_4700_) );
	OAI21X1 OAI21X1_315 ( .A(_3985_), .B(micro_hash_synth_2_W_21__6_), .C(_4630_), .Y(_4701_) );
	AOI21X1 AOI21X1_165 ( .A(_3985_), .B(micro_hash_synth_2_W_21__6_), .C(_4701_), .Y(_4702_) );
	OAI21X1 OAI21X1_316 ( .A(_4735__bF_buf9), .B(_4702_), .C(_4700_), .Y(_3200_) );
	NAND2X1 NAND2X1_183 ( .A(micro_hash_synth_2_W_30__7_), .B(_4269__bF_buf6), .Y(_4703_) );
	OAI21X1 OAI21X1_317 ( .A(_4452_), .B(micro_hash_synth_2_W_21__7_), .C(_4633_), .Y(_4704_) );
	AOI21X1 AOI21X1_166 ( .A(_4452_), .B(micro_hash_synth_2_W_21__7_), .C(_4704_), .Y(_4705_) );
	OAI21X1 OAI21X1_318 ( .A(_4735__bF_buf8), .B(_4705_), .C(_4703_), .Y(_3201_) );
	NAND2X1 NAND2X1_184 ( .A(micro_hash_synth_2_W_31__0_), .B(_4269__bF_buf5), .Y(_4706_) );
	OAI21X1 OAI21X1_319 ( .A(_4384_), .B(micro_hash_synth_2_W_22__0_), .C(_4636_), .Y(_4707_) );
	AOI21X1 AOI21X1_167 ( .A(_4384_), .B(micro_hash_synth_2_W_22__0_), .C(_4707_), .Y(_4708_) );
	OAI21X1 OAI21X1_320 ( .A(_4735__bF_buf7), .B(_4708_), .C(_4706_), .Y(_3202_) );
	OAI21X1 OAI21X1_321 ( .A(_4389_), .B(micro_hash_synth_2_W_22__1_), .C(_4639_), .Y(_4709_) );
	AOI21X1 AOI21X1_168 ( .A(_4389_), .B(micro_hash_synth_2_W_22__1_), .C(_4709_), .Y(_4710_) );
	OAI22X1 OAI22X1_206 ( .A(_4735__bF_buf6), .B(_4710_), .C(_4740__bF_buf0), .D(_3529_), .Y(_3203_) );
	OAI21X1 OAI21X1_322 ( .A(_4394_), .B(micro_hash_synth_2_W_22__2_), .C(_4642_), .Y(_4711_) );
	AOI21X1 AOI21X1_169 ( .A(_4394_), .B(micro_hash_synth_2_W_22__2_), .C(_4711_), .Y(_4712_) );
	OAI22X1 OAI22X1_207 ( .A(_4735__bF_buf5), .B(_4712_), .C(_4740__bF_buf13), .D(_3679_), .Y(_3204_) );
	NAND2X1 NAND2X1_185 ( .A(micro_hash_synth_2_W_31__3_), .B(_4269__bF_buf4), .Y(_4713_) );
	OAI21X1 OAI21X1_323 ( .A(_4399_), .B(micro_hash_synth_2_W_22__3_), .C(_4645_), .Y(_4714_) );
	AOI21X1 AOI21X1_170 ( .A(_4399_), .B(micro_hash_synth_2_W_22__3_), .C(_4714_), .Y(_4715_) );
	OAI21X1 OAI21X1_324 ( .A(_4735__bF_buf4), .B(_4715_), .C(_4713_), .Y(_3205_) );
	NAND2X1 NAND2X1_186 ( .A(micro_hash_synth_2_W_31__4_), .B(_4269__bF_buf3), .Y(_4716_) );
	OAI21X1 OAI21X1_325 ( .A(_4404_), .B(micro_hash_synth_2_W_22__4_), .C(_4648_), .Y(_4717_) );
	AOI21X1 AOI21X1_171 ( .A(_4404_), .B(micro_hash_synth_2_W_22__4_), .C(_4717_), .Y(_4718_) );
	OAI21X1 OAI21X1_326 ( .A(_4735__bF_buf3), .B(_4718_), .C(_4716_), .Y(_3206_) );
	NAND2X1 NAND2X1_187 ( .A(micro_hash_synth_2_W_31__5_), .B(_4269__bF_buf2), .Y(_4719_) );
	OAI21X1 OAI21X1_327 ( .A(_4409_), .B(micro_hash_synth_2_W_22__5_), .C(_4651_), .Y(_4720_) );
	AOI21X1 AOI21X1_172 ( .A(_4409_), .B(micro_hash_synth_2_W_22__5_), .C(_4720_), .Y(_4721_) );
	OAI21X1 OAI21X1_328 ( .A(_4735__bF_buf2), .B(_4721_), .C(_4719_), .Y(_3207_) );
	NAND2X1 NAND2X1_188 ( .A(micro_hash_synth_2_W_31__6_), .B(_4269__bF_buf1), .Y(_4722_) );
	OAI21X1 OAI21X1_329 ( .A(_4413_), .B(micro_hash_synth_2_W_22__6_), .C(_4654_), .Y(_4723_) );
	AOI21X1 AOI21X1_173 ( .A(_4413_), .B(micro_hash_synth_2_W_22__6_), .C(_4723_), .Y(_4724_) );
	OAI21X1 OAI21X1_330 ( .A(_4735__bF_buf1), .B(_4724_), .C(_4722_), .Y(_3208_) );
	NAND2X1 NAND2X1_189 ( .A(micro_hash_synth_2_W_31__7_), .B(_4269__bF_buf0), .Y(_4725_) );
	OAI21X1 OAI21X1_331 ( .A(_4417_), .B(micro_hash_synth_2_W_22__7_), .C(_4657_), .Y(_4726_) );
	AOI21X1 AOI21X1_174 ( .A(_4417_), .B(micro_hash_synth_2_W_22__7_), .C(_4726_), .Y(_4727_) );
	OAI21X1 OAI21X1_332 ( .A(_4735__bF_buf0), .B(_4727_), .C(_4725_), .Y(_3209_) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(clk_bF_buf113), .D(_3242_), .Q(micro_hash_synth_2_W_22__0_) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(clk_bF_buf112), .D(_3243_), .Q(micro_hash_synth_2_W_22__1_) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(clk_bF_buf111), .D(_3245_), .Q(micro_hash_synth_2_W_22__2_) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(clk_bF_buf110), .D(_3246_), .Q(micro_hash_synth_2_W_22__3_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(clk_bF_buf109), .D(_3247_), .Q(micro_hash_synth_2_W_22__4_) );
	DFFPOSX1 DFFPOSX1_6 ( .CLK(clk_bF_buf108), .D(_3248_), .Q(micro_hash_synth_2_W_22__5_) );
	DFFPOSX1 DFFPOSX1_7 ( .CLK(clk_bF_buf107), .D(_3249_), .Q(micro_hash_synth_2_W_22__6_) );
	DFFPOSX1 DFFPOSX1_8 ( .CLK(clk_bF_buf106), .D(_3250_), .Q(micro_hash_synth_2_W_22__7_) );
	DFFPOSX1 DFFPOSX1_9 ( .CLK(clk_bF_buf105), .D(_3077_), .Q(micro_hash_synth_2_W_0__0_) );
	DFFPOSX1 DFFPOSX1_10 ( .CLK(clk_bF_buf104), .D(_3078_), .Q(micro_hash_synth_2_W_0__1_) );
	DFFPOSX1 DFFPOSX1_11 ( .CLK(clk_bF_buf103), .D(_3080_), .Q(micro_hash_synth_2_W_0__2_) );
	DFFPOSX1 DFFPOSX1_12 ( .CLK(clk_bF_buf102), .D(_3081_), .Q(micro_hash_synth_2_W_0__3_) );
	DFFPOSX1 DFFPOSX1_13 ( .CLK(clk_bF_buf101), .D(_3082_), .Q(micro_hash_synth_2_W_0__4_) );
	DFFPOSX1 DFFPOSX1_14 ( .CLK(clk_bF_buf100), .D(_3083_), .Q(micro_hash_synth_2_W_0__5_) );
	DFFPOSX1 DFFPOSX1_15 ( .CLK(clk_bF_buf99), .D(_3084_), .Q(micro_hash_synth_2_W_0__6_) );
	DFFPOSX1 DFFPOSX1_16 ( .CLK(clk_bF_buf98), .D(_3085_), .Q(micro_hash_synth_2_W_0__7_) );
	DFFPOSX1 DFFPOSX1_17 ( .CLK(clk_bF_buf97), .D(_3298_), .Q(micro_hash_synth_2_W_19__0_) );
	DFFPOSX1 DFFPOSX1_18 ( .CLK(clk_bF_buf96), .D(_3299_), .Q(micro_hash_synth_2_W_19__1_) );
	DFFPOSX1 DFFPOSX1_19 ( .CLK(clk_bF_buf95), .D(_3300_), .Q(micro_hash_synth_2_W_19__2_) );
	DFFPOSX1 DFFPOSX1_20 ( .CLK(clk_bF_buf94), .D(_3301_), .Q(micro_hash_synth_2_W_19__3_) );
	DFFPOSX1 DFFPOSX1_21 ( .CLK(clk_bF_buf93), .D(_3303_), .Q(micro_hash_synth_2_W_19__4_) );
	DFFPOSX1 DFFPOSX1_22 ( .CLK(clk_bF_buf92), .D(_3304_), .Q(micro_hash_synth_2_W_19__5_) );
	DFFPOSX1 DFFPOSX1_23 ( .CLK(clk_bF_buf91), .D(_3305_), .Q(micro_hash_synth_2_W_19__6_) );
	DFFPOSX1 DFFPOSX1_24 ( .CLK(clk_bF_buf90), .D(_3306_), .Q(micro_hash_synth_2_W_19__7_) );
	DFFPOSX1 DFFPOSX1_25 ( .CLK(clk_bF_buf89), .D(_3278_), .Q(micro_hash_synth_2_W_20__0_) );
	DFFPOSX1 DFFPOSX1_26 ( .CLK(clk_bF_buf88), .D(_3279_), .Q(micro_hash_synth_2_W_20__1_) );
	DFFPOSX1 DFFPOSX1_27 ( .CLK(clk_bF_buf87), .D(_3280_), .Q(micro_hash_synth_2_W_20__2_) );
	DFFPOSX1 DFFPOSX1_28 ( .CLK(clk_bF_buf86), .D(_3281_), .Q(micro_hash_synth_2_W_20__3_) );
	DFFPOSX1 DFFPOSX1_29 ( .CLK(clk_bF_buf85), .D(_3282_), .Q(micro_hash_synth_2_W_20__4_) );
	DFFPOSX1 DFFPOSX1_30 ( .CLK(clk_bF_buf84), .D(_3283_), .Q(micro_hash_synth_2_W_20__5_) );
	DFFPOSX1 DFFPOSX1_31 ( .CLK(clk_bF_buf83), .D(_3284_), .Q(micro_hash_synth_2_W_20__6_) );
	DFFPOSX1 DFFPOSX1_32 ( .CLK(clk_bF_buf82), .D(_3285_), .Q(micro_hash_synth_2_W_20__7_) );
	DFFPOSX1 DFFPOSX1_33 ( .CLK(clk_bF_buf81), .D(_3269_), .Q(micro_hash_synth_2_W_21__0_) );
	DFFPOSX1 DFFPOSX1_34 ( .CLK(clk_bF_buf80), .D(_3270_), .Q(micro_hash_synth_2_W_21__1_) );
	DFFPOSX1 DFFPOSX1_35 ( .CLK(clk_bF_buf79), .D(_3271_), .Q(micro_hash_synth_2_W_21__2_) );
	DFFPOSX1 DFFPOSX1_36 ( .CLK(clk_bF_buf78), .D(_3272_), .Q(micro_hash_synth_2_W_21__3_) );
	DFFPOSX1 DFFPOSX1_37 ( .CLK(clk_bF_buf77), .D(_3273_), .Q(micro_hash_synth_2_W_21__4_) );
	DFFPOSX1 DFFPOSX1_38 ( .CLK(clk_bF_buf76), .D(_3274_), .Q(micro_hash_synth_2_W_21__5_) );
	DFFPOSX1 DFFPOSX1_39 ( .CLK(clk_bF_buf75), .D(_3275_), .Q(micro_hash_synth_2_W_21__6_) );
	DFFPOSX1 DFFPOSX1_40 ( .CLK(clk_bF_buf74), .D(_3276_), .Q(micro_hash_synth_2_W_21__7_) );
	DFFPOSX1 DFFPOSX1_41 ( .CLK(clk_bF_buf73), .D(_3047__0_), .Q(Hhash_synth2_0_) );
	DFFPOSX1 DFFPOSX1_42 ( .CLK(clk_bF_buf72), .D(_3047__1_), .Q(Hhash_synth2_1_) );
	DFFPOSX1 DFFPOSX1_43 ( .CLK(clk_bF_buf71), .D(_3047__2_), .Q(Hhash_synth2_2_) );
	DFFPOSX1 DFFPOSX1_44 ( .CLK(clk_bF_buf70), .D(_3047__3_), .Q(Hhash_synth2_3_) );
	DFFPOSX1 DFFPOSX1_45 ( .CLK(clk_bF_buf69), .D(_3047__4_), .Q(Hhash_synth2_4_) );
	DFFPOSX1 DFFPOSX1_46 ( .CLK(clk_bF_buf68), .D(_3047__5_), .Q(Hhash_synth2_5_) );
	DFFPOSX1 DFFPOSX1_47 ( .CLK(clk_bF_buf67), .D(_3047__6_), .Q(Hhash_synth2_6_) );
	DFFPOSX1 DFFPOSX1_48 ( .CLK(clk_bF_buf66), .D(_3047__7_), .Q(Hhash_synth2_7_) );
	DFFPOSX1 DFFPOSX1_49 ( .CLK(clk_bF_buf65), .D(_3047__8_), .Q(Hhash_synth2_8_) );
	DFFPOSX1 DFFPOSX1_50 ( .CLK(clk_bF_buf64), .D(_3047__9_), .Q(Hhash_synth2_9_) );
	DFFPOSX1 DFFPOSX1_51 ( .CLK(clk_bF_buf63), .D(_3047__10_), .Q(Hhash_synth2_10_) );
	DFFPOSX1 DFFPOSX1_52 ( .CLK(clk_bF_buf62), .D(_3047__11_), .Q(Hhash_synth2_11_) );
	DFFPOSX1 DFFPOSX1_53 ( .CLK(clk_bF_buf61), .D(_3047__12_), .Q(Hhash_synth2_12_) );
	DFFPOSX1 DFFPOSX1_54 ( .CLK(clk_bF_buf60), .D(_3047__13_), .Q(Hhash_synth2_13_) );
	DFFPOSX1 DFFPOSX1_55 ( .CLK(clk_bF_buf59), .D(_3047__14_), .Q(Hhash_synth2_14_) );
	DFFPOSX1 DFFPOSX1_56 ( .CLK(clk_bF_buf58), .D(_3047__15_), .Q(Hhash_synth2_15_) );
	DFFPOSX1 DFFPOSX1_57 ( .CLK(clk_bF_buf57), .D(_3047__16_), .Q(Hhash_synth2_16_) );
	DFFPOSX1 DFFPOSX1_58 ( .CLK(clk_bF_buf56), .D(_3047__17_), .Q(Hhash_synth2_17_) );
	DFFPOSX1 DFFPOSX1_59 ( .CLK(clk_bF_buf55), .D(_3047__18_), .Q(Hhash_synth2_18_) );
	DFFPOSX1 DFFPOSX1_60 ( .CLK(clk_bF_buf54), .D(_3047__19_), .Q(Hhash_synth2_19_) );
	DFFPOSX1 DFFPOSX1_61 ( .CLK(clk_bF_buf53), .D(_3047__20_), .Q(Hhash_synth2_20_) );
	DFFPOSX1 DFFPOSX1_62 ( .CLK(clk_bF_buf52), .D(_3047__21_), .Q(Hhash_synth2_21_) );
	DFFPOSX1 DFFPOSX1_63 ( .CLK(clk_bF_buf51), .D(_3047__22_), .Q(Hhash_synth2_22_) );
	DFFPOSX1 DFFPOSX1_64 ( .CLK(clk_bF_buf50), .D(_3047__23_), .Q(Hhash_synth2_23_) );
	DFFPOSX1 DFFPOSX1_65 ( .CLK(clk_bF_buf49), .D(_3052__0_), .Q(micro_hash_synth_2_nonce_synth_1_0_) );
	DFFPOSX1 DFFPOSX1_66 ( .CLK(clk_bF_buf48), .D(_3052__1_), .Q(micro_hash_synth_2_nonce_synth_1_1_) );
	DFFPOSX1 DFFPOSX1_67 ( .CLK(clk_bF_buf47), .D(_3052__2_), .Q(micro_hash_synth_2_nonce_synth_1_2_) );
	DFFPOSX1 DFFPOSX1_68 ( .CLK(clk_bF_buf46), .D(_3052__3_), .Q(micro_hash_synth_2_nonce_synth_1_3_) );
	DFFPOSX1 DFFPOSX1_69 ( .CLK(clk_bF_buf45), .D(_3052__4_), .Q(micro_hash_synth_2_nonce_synth_1_4_) );
	DFFPOSX1 DFFPOSX1_70 ( .CLK(clk_bF_buf44), .D(_3052__5_), .Q(micro_hash_synth_2_nonce_synth_1_5_) );
	DFFPOSX1 DFFPOSX1_71 ( .CLK(clk_bF_buf43), .D(_3052__6_), .Q(micro_hash_synth_2_nonce_synth_1_6_) );
	DFFPOSX1 DFFPOSX1_72 ( .CLK(clk_bF_buf42), .D(_3052__7_), .Q(micro_hash_synth_2_nonce_synth_1_7_) );
	DFFPOSX1 DFFPOSX1_73 ( .CLK(clk_bF_buf41), .D(_3052__8_), .Q(micro_hash_synth_2_nonce_synth_1_8_) );
	DFFPOSX1 DFFPOSX1_74 ( .CLK(clk_bF_buf40), .D(_3052__9_), .Q(micro_hash_synth_2_nonce_synth_1_9_) );
	DFFPOSX1 DFFPOSX1_75 ( .CLK(clk_bF_buf39), .D(_3052__10_), .Q(micro_hash_synth_2_nonce_synth_1_10_) );
	DFFPOSX1 DFFPOSX1_76 ( .CLK(clk_bF_buf38), .D(_3052__11_), .Q(micro_hash_synth_2_nonce_synth_1_11_) );
	DFFPOSX1 DFFPOSX1_77 ( .CLK(clk_bF_buf37), .D(_3052__12_), .Q(micro_hash_synth_2_nonce_synth_1_12_) );
	DFFPOSX1 DFFPOSX1_78 ( .CLK(clk_bF_buf36), .D(_3052__13_), .Q(micro_hash_synth_2_nonce_synth_1_13_) );
	DFFPOSX1 DFFPOSX1_79 ( .CLK(clk_bF_buf35), .D(_3052__14_), .Q(micro_hash_synth_2_nonce_synth_1_14_) );
	DFFPOSX1 DFFPOSX1_80 ( .CLK(clk_bF_buf34), .D(_3052__15_), .Q(micro_hash_synth_2_nonce_synth_1_15_) );
	DFFPOSX1 DFFPOSX1_81 ( .CLK(clk_bF_buf33), .D(_3052__16_), .Q(micro_hash_synth_2_nonce_synth_1_16_) );
	DFFPOSX1 DFFPOSX1_82 ( .CLK(clk_bF_buf32), .D(_3052__17_), .Q(micro_hash_synth_2_nonce_synth_1_17_) );
	DFFPOSX1 DFFPOSX1_83 ( .CLK(clk_bF_buf31), .D(_3052__18_), .Q(micro_hash_synth_2_nonce_synth_1_18_) );
	DFFPOSX1 DFFPOSX1_84 ( .CLK(clk_bF_buf30), .D(_3052__19_), .Q(micro_hash_synth_2_nonce_synth_1_19_) );
	DFFPOSX1 DFFPOSX1_85 ( .CLK(clk_bF_buf29), .D(_3052__20_), .Q(micro_hash_synth_2_nonce_synth_1_20_) );
	DFFPOSX1 DFFPOSX1_86 ( .CLK(clk_bF_buf28), .D(_3052__21_), .Q(micro_hash_synth_2_nonce_synth_1_21_) );
	DFFPOSX1 DFFPOSX1_87 ( .CLK(clk_bF_buf27), .D(_3052__22_), .Q(micro_hash_synth_2_nonce_synth_1_22_) );
	DFFPOSX1 DFFPOSX1_88 ( .CLK(clk_bF_buf26), .D(_3052__23_), .Q(micro_hash_synth_2_nonce_synth_1_23_) );
	DFFPOSX1 DFFPOSX1_89 ( .CLK(clk_bF_buf25), .D(_3052__24_), .Q(micro_hash_synth_2_nonce_synth_1_24_) );
	DFFPOSX1 DFFPOSX1_90 ( .CLK(clk_bF_buf24), .D(_3052__25_), .Q(micro_hash_synth_2_nonce_synth_1_25_) );
	DFFPOSX1 DFFPOSX1_91 ( .CLK(clk_bF_buf23), .D(_3052__26_), .Q(micro_hash_synth_2_nonce_synth_1_26_) );
	DFFPOSX1 DFFPOSX1_92 ( .CLK(clk_bF_buf22), .D(_3052__27_), .Q(micro_hash_synth_2_nonce_synth_1_27_) );
	DFFPOSX1 DFFPOSX1_93 ( .CLK(clk_bF_buf21), .D(_3052__28_), .Q(micro_hash_synth_2_nonce_synth_1_28_) );
	DFFPOSX1 DFFPOSX1_94 ( .CLK(clk_bF_buf20), .D(_3052__29_), .Q(micro_hash_synth_2_nonce_synth_1_29_) );
	DFFPOSX1 DFFPOSX1_95 ( .CLK(clk_bF_buf19), .D(_3052__30_), .Q(micro_hash_synth_2_nonce_synth_1_30_) );
	DFFPOSX1 DFFPOSX1_96 ( .CLK(clk_bF_buf18), .D(_3052__31_), .Q(micro_hash_synth_2_nonce_synth_1_31_) );
	DFFPOSX1 DFFPOSX1_97 ( .CLK(clk_bF_buf17), .D(_3048__0_), .Q(micro_hash_synth_2_a_0_) );
	DFFPOSX1 DFFPOSX1_98 ( .CLK(clk_bF_buf16), .D(_3048__1_), .Q(micro_hash_synth_2_a_1_) );
	DFFPOSX1 DFFPOSX1_99 ( .CLK(clk_bF_buf15), .D(_3048__2_), .Q(micro_hash_synth_2_a_2_) );
	DFFPOSX1 DFFPOSX1_100 ( .CLK(clk_bF_buf14), .D(_3048__3_), .Q(micro_hash_synth_2_a_3_) );
	DFFPOSX1 DFFPOSX1_101 ( .CLK(clk_bF_buf13), .D(_3048__4_), .Q(micro_hash_synth_2_a_4_) );
	DFFPOSX1 DFFPOSX1_102 ( .CLK(clk_bF_buf12), .D(_3048__5_), .Q(micro_hash_synth_2_a_5_) );
	DFFPOSX1 DFFPOSX1_103 ( .CLK(clk_bF_buf11), .D(_3048__6_), .Q(micro_hash_synth_2_a_6_) );
	DFFPOSX1 DFFPOSX1_104 ( .CLK(clk_bF_buf10), .D(_3048__7_), .Q(micro_hash_synth_2_a_7_) );
	DFFPOSX1 DFFPOSX1_105 ( .CLK(clk_bF_buf9), .D(_3049__0_), .Q(micro_hash_synth_2_b_0_) );
	DFFPOSX1 DFFPOSX1_106 ( .CLK(clk_bF_buf8), .D(_3049__1_), .Q(micro_hash_synth_2_b_1_) );
	DFFPOSX1 DFFPOSX1_107 ( .CLK(clk_bF_buf7), .D(_3049__2_), .Q(micro_hash_synth_2_b_2_) );
	DFFPOSX1 DFFPOSX1_108 ( .CLK(clk_bF_buf6), .D(_3049__3_), .Q(micro_hash_synth_2_b_3_) );
	DFFPOSX1 DFFPOSX1_109 ( .CLK(clk_bF_buf5), .D(_3049__4_), .Q(micro_hash_synth_2_b_4_) );
	DFFPOSX1 DFFPOSX1_110 ( .CLK(clk_bF_buf4), .D(_3049__5_), .Q(micro_hash_synth_2_b_5_) );
	DFFPOSX1 DFFPOSX1_111 ( .CLK(clk_bF_buf3), .D(_3049__6_), .Q(micro_hash_synth_2_b_6_) );
	DFFPOSX1 DFFPOSX1_112 ( .CLK(clk_bF_buf2), .D(_3049__7_), .Q(micro_hash_synth_2_b_7_) );
	DFFPOSX1 DFFPOSX1_113 ( .CLK(clk_bF_buf1), .D(_3050__0_), .Q(micro_hash_synth_2_c_0_) );
	DFFPOSX1 DFFPOSX1_114 ( .CLK(clk_bF_buf0), .D(_3050__1_), .Q(micro_hash_synth_2_c_1_) );
	DFFPOSX1 DFFPOSX1_115 ( .CLK(clk_bF_buf113), .D(_3050__2_), .Q(micro_hash_synth_2_c_2_) );
	DFFPOSX1 DFFPOSX1_116 ( .CLK(clk_bF_buf112), .D(_3050__3_), .Q(micro_hash_synth_2_c_3_) );
	DFFPOSX1 DFFPOSX1_117 ( .CLK(clk_bF_buf111), .D(_3050__4_), .Q(micro_hash_synth_2_c_4_) );
	DFFPOSX1 DFFPOSX1_118 ( .CLK(clk_bF_buf110), .D(_3050__5_), .Q(micro_hash_synth_2_c_5_) );
	DFFPOSX1 DFFPOSX1_119 ( .CLK(clk_bF_buf109), .D(_3050__6_), .Q(micro_hash_synth_2_c_6_) );
	DFFPOSX1 DFFPOSX1_120 ( .CLK(clk_bF_buf108), .D(_3050__7_), .Q(micro_hash_synth_2_c_7_) );
	DFFPOSX1 DFFPOSX1_121 ( .CLK(clk_bF_buf107), .D(_3051__0_), .Q(micro_hash_synth_2_k_0_) );
	DFFPOSX1 DFFPOSX1_122 ( .CLK(clk_bF_buf106), .D(_3051__1_), .Q(micro_hash_synth_2_k_1_) );
	DFFPOSX1 DFFPOSX1_123 ( .CLK(clk_bF_buf105), .D(_3051__2_), .Q(micro_hash_synth_2_k_2_) );
	DFFPOSX1 DFFPOSX1_124 ( .CLK(clk_bF_buf104), .D(_3051__3_), .Q(micro_hash_synth_2_k_3_) );
	DFFPOSX1 DFFPOSX1_125 ( .CLK(clk_bF_buf103), .D(_3051__4_), .Q(micro_hash_synth_2_k_4_) );
	DFFPOSX1 DFFPOSX1_126 ( .CLK(clk_bF_buf102), .D(_3051__5_), .Q(micro_hash_synth_2_k_5_) );
	DFFPOSX1 DFFPOSX1_127 ( .CLK(clk_bF_buf101), .D(_3051__6_), .Q(micro_hash_synth_2_k_6_) );
	DFFPOSX1 DFFPOSX1_128 ( .CLK(clk_bF_buf100), .D(_3051__7_), .Q(micro_hash_synth_2_k_7_) );
	DFFPOSX1 DFFPOSX1_129 ( .CLK(clk_bF_buf99), .D(_3053__0_), .Q(micro_hash_synth_2_x_0_) );
	DFFPOSX1 DFFPOSX1_130 ( .CLK(clk_bF_buf98), .D(_3053__1_), .Q(micro_hash_synth_2_x_1_) );
	DFFPOSX1 DFFPOSX1_131 ( .CLK(clk_bF_buf97), .D(_3053__2_), .Q(micro_hash_synth_2_x_2_) );
	DFFPOSX1 DFFPOSX1_132 ( .CLK(clk_bF_buf96), .D(_3053__3_), .Q(micro_hash_synth_2_x_3_) );
	DFFPOSX1 DFFPOSX1_133 ( .CLK(clk_bF_buf95), .D(_3053__4_), .Q(micro_hash_synth_2_x_4_) );
	DFFPOSX1 DFFPOSX1_134 ( .CLK(clk_bF_buf94), .D(_3053__5_), .Q(micro_hash_synth_2_x_5_) );
	DFFPOSX1 DFFPOSX1_135 ( .CLK(clk_bF_buf93), .D(_3053__6_), .Q(micro_hash_synth_2_x_6_) );
	DFFPOSX1 DFFPOSX1_136 ( .CLK(clk_bF_buf92), .D(_3053__7_), .Q(micro_hash_synth_2_x_7_) );
	DFFPOSX1 DFFPOSX1_137 ( .CLK(clk_bF_buf91), .D(_3086_), .Q(micro_hash_synth_2_W_18__0_) );
	DFFPOSX1 DFFPOSX1_138 ( .CLK(clk_bF_buf90), .D(_3087_), .Q(micro_hash_synth_2_W_18__1_) );
	DFFPOSX1 DFFPOSX1_139 ( .CLK(clk_bF_buf89), .D(_3088_), .Q(micro_hash_synth_2_W_18__2_) );
	DFFPOSX1 DFFPOSX1_140 ( .CLK(clk_bF_buf88), .D(_3089_), .Q(micro_hash_synth_2_W_18__3_) );
	DFFPOSX1 DFFPOSX1_141 ( .CLK(clk_bF_buf87), .D(_3090_), .Q(micro_hash_synth_2_W_18__4_) );
	DFFPOSX1 DFFPOSX1_142 ( .CLK(clk_bF_buf86), .D(_3091_), .Q(micro_hash_synth_2_W_18__5_) );
	DFFPOSX1 DFFPOSX1_143 ( .CLK(clk_bF_buf85), .D(_3092_), .Q(micro_hash_synth_2_W_18__6_) );
	DFFPOSX1 DFFPOSX1_144 ( .CLK(clk_bF_buf84), .D(_3093_), .Q(micro_hash_synth_2_W_18__7_) );
	DFFPOSX1 DFFPOSX1_145 ( .CLK(clk_bF_buf83), .D(_3094_), .Q(micro_hash_synth_2_W_17__0_) );
	DFFPOSX1 DFFPOSX1_146 ( .CLK(clk_bF_buf82), .D(_3096_), .Q(micro_hash_synth_2_W_17__1_) );
	DFFPOSX1 DFFPOSX1_147 ( .CLK(clk_bF_buf81), .D(_3097_), .Q(micro_hash_synth_2_W_17__2_) );
	DFFPOSX1 DFFPOSX1_148 ( .CLK(clk_bF_buf80), .D(_3098_), .Q(micro_hash_synth_2_W_17__3_) );
	DFFPOSX1 DFFPOSX1_149 ( .CLK(clk_bF_buf79), .D(_3099_), .Q(micro_hash_synth_2_W_17__4_) );
	DFFPOSX1 DFFPOSX1_150 ( .CLK(clk_bF_buf78), .D(_3100_), .Q(micro_hash_synth_2_W_17__5_) );
	DFFPOSX1 DFFPOSX1_151 ( .CLK(clk_bF_buf77), .D(_3101_), .Q(micro_hash_synth_2_W_17__6_) );
	DFFPOSX1 DFFPOSX1_152 ( .CLK(clk_bF_buf76), .D(_3102_), .Q(micro_hash_synth_2_W_17__7_) );
	DFFPOSX1 DFFPOSX1_153 ( .CLK(clk_bF_buf75), .D(_3129_), .Q(micro_hash_synth_2_W_16__0_) );
	DFFPOSX1 DFFPOSX1_154 ( .CLK(clk_bF_buf74), .D(_3130_), .Q(micro_hash_synth_2_W_16__1_) );
	DFFPOSX1 DFFPOSX1_155 ( .CLK(clk_bF_buf73), .D(_3131_), .Q(micro_hash_synth_2_W_16__2_) );
	DFFPOSX1 DFFPOSX1_156 ( .CLK(clk_bF_buf72), .D(_3132_), .Q(micro_hash_synth_2_W_16__3_) );
	DFFPOSX1 DFFPOSX1_157 ( .CLK(clk_bF_buf71), .D(_3133_), .Q(micro_hash_synth_2_W_16__4_) );
	DFFPOSX1 DFFPOSX1_158 ( .CLK(clk_bF_buf70), .D(_3134_), .Q(micro_hash_synth_2_W_16__5_) );
	DFFPOSX1 DFFPOSX1_159 ( .CLK(clk_bF_buf69), .D(_3135_), .Q(micro_hash_synth_2_W_16__6_) );
	DFFPOSX1 DFFPOSX1_160 ( .CLK(clk_bF_buf68), .D(_3136_), .Q(micro_hash_synth_2_W_16__7_) );
	DFFPOSX1 DFFPOSX1_161 ( .CLK(clk_bF_buf67), .D(_3103_), .Q(micro_hash_synth_2_W_15__0_) );
	DFFPOSX1 DFFPOSX1_162 ( .CLK(clk_bF_buf66), .D(_3104_), .Q(micro_hash_synth_2_W_15__1_) );
	DFFPOSX1 DFFPOSX1_163 ( .CLK(clk_bF_buf65), .D(_3105_), .Q(micro_hash_synth_2_W_15__2_) );
	DFFPOSX1 DFFPOSX1_164 ( .CLK(clk_bF_buf64), .D(_3106_), .Q(micro_hash_synth_2_W_15__3_) );
	DFFPOSX1 DFFPOSX1_165 ( .CLK(clk_bF_buf63), .D(_3107_), .Q(micro_hash_synth_2_W_15__4_) );
	DFFPOSX1 DFFPOSX1_166 ( .CLK(clk_bF_buf62), .D(_3108_), .Q(micro_hash_synth_2_W_15__5_) );
	DFFPOSX1 DFFPOSX1_167 ( .CLK(clk_bF_buf61), .D(_3109_), .Q(micro_hash_synth_2_W_15__6_) );
	DFFPOSX1 DFFPOSX1_168 ( .CLK(clk_bF_buf60), .D(_3110_), .Q(micro_hash_synth_2_W_15__7_) );
	DFFPOSX1 DFFPOSX1_169 ( .CLK(clk_bF_buf59), .D(_3068_), .Q(micro_hash_synth_2_W_14__0_) );
	DFFPOSX1 DFFPOSX1_170 ( .CLK(clk_bF_buf58), .D(_3069_), .Q(micro_hash_synth_2_W_14__1_) );
	DFFPOSX1 DFFPOSX1_171 ( .CLK(clk_bF_buf57), .D(_3070_), .Q(micro_hash_synth_2_W_14__2_) );
	DFFPOSX1 DFFPOSX1_172 ( .CLK(clk_bF_buf56), .D(_3071_), .Q(micro_hash_synth_2_W_14__3_) );
	DFFPOSX1 DFFPOSX1_173 ( .CLK(clk_bF_buf55), .D(_3072_), .Q(micro_hash_synth_2_W_14__4_) );
	DFFPOSX1 DFFPOSX1_174 ( .CLK(clk_bF_buf54), .D(_3073_), .Q(micro_hash_synth_2_W_14__5_) );
	DFFPOSX1 DFFPOSX1_175 ( .CLK(clk_bF_buf53), .D(_3074_), .Q(micro_hash_synth_2_W_14__6_) );
	DFFPOSX1 DFFPOSX1_176 ( .CLK(clk_bF_buf52), .D(_3075_), .Q(micro_hash_synth_2_W_14__7_) );
	DFFPOSX1 DFFPOSX1_177 ( .CLK(clk_bF_buf51), .D(_3120_), .Q(micro_hash_synth_2_W_13__0_) );
	DFFPOSX1 DFFPOSX1_178 ( .CLK(clk_bF_buf50), .D(_3121_), .Q(micro_hash_synth_2_W_13__1_) );
	DFFPOSX1 DFFPOSX1_179 ( .CLK(clk_bF_buf49), .D(_3122_), .Q(micro_hash_synth_2_W_13__2_) );
	DFFPOSX1 DFFPOSX1_180 ( .CLK(clk_bF_buf48), .D(_3123_), .Q(micro_hash_synth_2_W_13__3_) );
	DFFPOSX1 DFFPOSX1_181 ( .CLK(clk_bF_buf47), .D(_3124_), .Q(micro_hash_synth_2_W_13__4_) );
	DFFPOSX1 DFFPOSX1_182 ( .CLK(clk_bF_buf46), .D(_3125_), .Q(micro_hash_synth_2_W_13__5_) );
	DFFPOSX1 DFFPOSX1_183 ( .CLK(clk_bF_buf45), .D(_3126_), .Q(micro_hash_synth_2_W_13__6_) );
	DFFPOSX1 DFFPOSX1_184 ( .CLK(clk_bF_buf44), .D(_3128_), .Q(micro_hash_synth_2_W_13__7_) );
	DFFPOSX1 DFFPOSX1_185 ( .CLK(clk_bF_buf43), .D(_3286_), .Q(micro_hash_synth_2_W_12__0_) );
	DFFPOSX1 DFFPOSX1_186 ( .CLK(clk_bF_buf42), .D(_3287_), .Q(micro_hash_synth_2_W_12__1_) );
	DFFPOSX1 DFFPOSX1_187 ( .CLK(clk_bF_buf41), .D(_3289_), .Q(micro_hash_synth_2_W_12__2_) );
	DFFPOSX1 DFFPOSX1_188 ( .CLK(clk_bF_buf40), .D(_3290_), .Q(micro_hash_synth_2_W_12__3_) );
	DFFPOSX1 DFFPOSX1_189 ( .CLK(clk_bF_buf39), .D(_3291_), .Q(micro_hash_synth_2_W_12__4_) );
	DFFPOSX1 DFFPOSX1_190 ( .CLK(clk_bF_buf38), .D(_3292_), .Q(micro_hash_synth_2_W_12__5_) );
	DFFPOSX1 DFFPOSX1_191 ( .CLK(clk_bF_buf37), .D(_3293_), .Q(micro_hash_synth_2_W_12__6_) );
	DFFPOSX1 DFFPOSX1_192 ( .CLK(clk_bF_buf36), .D(_3294_), .Q(micro_hash_synth_2_W_12__7_) );
	DFFPOSX1 DFFPOSX1_193 ( .CLK(clk_bF_buf35), .D(_3154_), .Q(micro_hash_synth_2_W_11__0_) );
	DFFPOSX1 DFFPOSX1_194 ( .CLK(clk_bF_buf34), .D(_3155_), .Q(micro_hash_synth_2_W_11__1_) );
	DFFPOSX1 DFFPOSX1_195 ( .CLK(clk_bF_buf33), .D(_3156_), .Q(micro_hash_synth_2_W_11__2_) );
	DFFPOSX1 DFFPOSX1_196 ( .CLK(clk_bF_buf32), .D(_3157_), .Q(micro_hash_synth_2_W_11__3_) );
	DFFPOSX1 DFFPOSX1_197 ( .CLK(clk_bF_buf31), .D(_3158_), .Q(micro_hash_synth_2_W_11__4_) );
	DFFPOSX1 DFFPOSX1_198 ( .CLK(clk_bF_buf30), .D(_3159_), .Q(micro_hash_synth_2_W_11__5_) );
	DFFPOSX1 DFFPOSX1_199 ( .CLK(clk_bF_buf29), .D(_3160_), .Q(micro_hash_synth_2_W_11__6_) );
	DFFPOSX1 DFFPOSX1_200 ( .CLK(clk_bF_buf28), .D(_3161_), .Q(micro_hash_synth_2_W_11__7_) );
	DFFPOSX1 DFFPOSX1_201 ( .CLK(clk_bF_buf27), .D(_3146_), .Q(micro_hash_synth_2_W_10__0_) );
	DFFPOSX1 DFFPOSX1_202 ( .CLK(clk_bF_buf26), .D(_3147_), .Q(micro_hash_synth_2_W_10__1_) );
	DFFPOSX1 DFFPOSX1_203 ( .CLK(clk_bF_buf25), .D(_3148_), .Q(micro_hash_synth_2_W_10__2_) );
	DFFPOSX1 DFFPOSX1_204 ( .CLK(clk_bF_buf24), .D(_3149_), .Q(micro_hash_synth_2_W_10__3_) );
	DFFPOSX1 DFFPOSX1_205 ( .CLK(clk_bF_buf23), .D(_3150_), .Q(micro_hash_synth_2_W_10__4_) );
	DFFPOSX1 DFFPOSX1_206 ( .CLK(clk_bF_buf22), .D(_3151_), .Q(micro_hash_synth_2_W_10__5_) );
	DFFPOSX1 DFFPOSX1_207 ( .CLK(clk_bF_buf21), .D(_3152_), .Q(micro_hash_synth_2_W_10__6_) );
	DFFPOSX1 DFFPOSX1_208 ( .CLK(clk_bF_buf20), .D(_3153_), .Q(micro_hash_synth_2_W_10__7_) );
	DFFPOSX1 DFFPOSX1_209 ( .CLK(clk_bF_buf19), .D(_3251_), .Q(micro_hash_synth_2_W_9__0_) );
	DFFPOSX1 DFFPOSX1_210 ( .CLK(clk_bF_buf18), .D(_3252_), .Q(micro_hash_synth_2_W_9__1_) );
	DFFPOSX1 DFFPOSX1_211 ( .CLK(clk_bF_buf17), .D(_3253_), .Q(micro_hash_synth_2_W_9__2_) );
	DFFPOSX1 DFFPOSX1_212 ( .CLK(clk_bF_buf16), .D(_3254_), .Q(micro_hash_synth_2_W_9__3_) );
	DFFPOSX1 DFFPOSX1_213 ( .CLK(clk_bF_buf15), .D(_3256_), .Q(micro_hash_synth_2_W_9__4_) );
	DFFPOSX1 DFFPOSX1_214 ( .CLK(clk_bF_buf14), .D(_3257_), .Q(micro_hash_synth_2_W_9__5_) );
	DFFPOSX1 DFFPOSX1_215 ( .CLK(clk_bF_buf13), .D(_3258_), .Q(micro_hash_synth_2_W_9__6_) );
	DFFPOSX1 DFFPOSX1_216 ( .CLK(clk_bF_buf12), .D(_3259_), .Q(micro_hash_synth_2_W_9__7_) );
	DFFPOSX1 DFFPOSX1_217 ( .CLK(clk_bF_buf11), .D(_3302_), .Q(micro_hash_synth_2_W_8__0_) );
	DFFPOSX1 DFFPOSX1_218 ( .CLK(clk_bF_buf10), .D(_3307_), .Q(micro_hash_synth_2_W_8__1_) );
	DFFPOSX1 DFFPOSX1_219 ( .CLK(clk_bF_buf9), .D(_3308_), .Q(micro_hash_synth_2_W_8__2_) );
	DFFPOSX1 DFFPOSX1_220 ( .CLK(clk_bF_buf8), .D(_3309_), .Q(micro_hash_synth_2_W_8__3_) );
	DFFPOSX1 DFFPOSX1_221 ( .CLK(clk_bF_buf7), .D(_3054_), .Q(micro_hash_synth_2_W_8__4_) );
	DFFPOSX1 DFFPOSX1_222 ( .CLK(clk_bF_buf6), .D(_3055_), .Q(micro_hash_synth_2_W_8__5_) );
	DFFPOSX1 DFFPOSX1_223 ( .CLK(clk_bF_buf5), .D(_3063_), .Q(micro_hash_synth_2_W_8__6_) );
	DFFPOSX1 DFFPOSX1_224 ( .CLK(clk_bF_buf4), .D(_3065_), .Q(micro_hash_synth_2_W_8__7_) );
	DFFPOSX1 DFFPOSX1_225 ( .CLK(clk_bF_buf3), .D(_3234_), .Q(micro_hash_synth_2_W_7__0_) );
	DFFPOSX1 DFFPOSX1_226 ( .CLK(clk_bF_buf2), .D(_3235_), .Q(micro_hash_synth_2_W_7__1_) );
	DFFPOSX1 DFFPOSX1_227 ( .CLK(clk_bF_buf1), .D(_3236_), .Q(micro_hash_synth_2_W_7__2_) );
	DFFPOSX1 DFFPOSX1_228 ( .CLK(clk_bF_buf0), .D(_3237_), .Q(micro_hash_synth_2_W_7__3_) );
	DFFPOSX1 DFFPOSX1_229 ( .CLK(clk_bF_buf113), .D(_3238_), .Q(micro_hash_synth_2_W_7__4_) );
	DFFPOSX1 DFFPOSX1_230 ( .CLK(clk_bF_buf112), .D(_3239_), .Q(micro_hash_synth_2_W_7__5_) );
	DFFPOSX1 DFFPOSX1_231 ( .CLK(clk_bF_buf111), .D(_3240_), .Q(micro_hash_synth_2_W_7__6_) );
	DFFPOSX1 DFFPOSX1_232 ( .CLK(clk_bF_buf110), .D(_3241_), .Q(micro_hash_synth_2_W_7__7_) );
	DFFPOSX1 DFFPOSX1_233 ( .CLK(clk_bF_buf109), .D(_3112_), .Q(micro_hash_synth_2_W_6__0_) );
	DFFPOSX1 DFFPOSX1_234 ( .CLK(clk_bF_buf108), .D(_3113_), .Q(micro_hash_synth_2_W_6__1_) );
	DFFPOSX1 DFFPOSX1_235 ( .CLK(clk_bF_buf107), .D(_3114_), .Q(micro_hash_synth_2_W_6__2_) );
	DFFPOSX1 DFFPOSX1_236 ( .CLK(clk_bF_buf106), .D(_3115_), .Q(micro_hash_synth_2_W_6__3_) );
	DFFPOSX1 DFFPOSX1_237 ( .CLK(clk_bF_buf105), .D(_3116_), .Q(micro_hash_synth_2_W_6__4_) );
	DFFPOSX1 DFFPOSX1_238 ( .CLK(clk_bF_buf104), .D(_3117_), .Q(micro_hash_synth_2_W_6__5_) );
	DFFPOSX1 DFFPOSX1_239 ( .CLK(clk_bF_buf103), .D(_3118_), .Q(micro_hash_synth_2_W_6__6_) );
	DFFPOSX1 DFFPOSX1_240 ( .CLK(clk_bF_buf102), .D(_3119_), .Q(micro_hash_synth_2_W_6__7_) );
	DFFPOSX1 DFFPOSX1_241 ( .CLK(clk_bF_buf101), .D(_3056_), .Q(micro_hash_synth_2_W_5__0_) );
	DFFPOSX1 DFFPOSX1_242 ( .CLK(clk_bF_buf100), .D(_3057_), .Q(micro_hash_synth_2_W_5__1_) );
	DFFPOSX1 DFFPOSX1_243 ( .CLK(clk_bF_buf99), .D(_3058_), .Q(micro_hash_synth_2_W_5__2_) );
	DFFPOSX1 DFFPOSX1_244 ( .CLK(clk_bF_buf98), .D(_3059_), .Q(micro_hash_synth_2_W_5__3_) );
	DFFPOSX1 DFFPOSX1_245 ( .CLK(clk_bF_buf97), .D(_3060_), .Q(micro_hash_synth_2_W_5__4_) );
	DFFPOSX1 DFFPOSX1_246 ( .CLK(clk_bF_buf96), .D(_3061_), .Q(micro_hash_synth_2_W_5__5_) );
	DFFPOSX1 DFFPOSX1_247 ( .CLK(clk_bF_buf95), .D(_3062_), .Q(micro_hash_synth_2_W_5__6_) );
	DFFPOSX1 DFFPOSX1_248 ( .CLK(clk_bF_buf94), .D(_3064_), .Q(micro_hash_synth_2_W_5__7_) );
	DFFPOSX1 DFFPOSX1_249 ( .CLK(clk_bF_buf93), .D(_3260_), .Q(micro_hash_synth_2_W_4__0_) );
	DFFPOSX1 DFFPOSX1_250 ( .CLK(clk_bF_buf92), .D(_3261_), .Q(micro_hash_synth_2_W_4__1_) );
	DFFPOSX1 DFFPOSX1_251 ( .CLK(clk_bF_buf91), .D(_3262_), .Q(micro_hash_synth_2_W_4__2_) );
	DFFPOSX1 DFFPOSX1_252 ( .CLK(clk_bF_buf90), .D(_3263_), .Q(micro_hash_synth_2_W_4__3_) );
	DFFPOSX1 DFFPOSX1_253 ( .CLK(clk_bF_buf89), .D(_3264_), .Q(micro_hash_synth_2_W_4__4_) );
	DFFPOSX1 DFFPOSX1_254 ( .CLK(clk_bF_buf88), .D(_3265_), .Q(micro_hash_synth_2_W_4__5_) );
	DFFPOSX1 DFFPOSX1_255 ( .CLK(clk_bF_buf87), .D(_3267_), .Q(micro_hash_synth_2_W_4__6_) );
	DFFPOSX1 DFFPOSX1_256 ( .CLK(clk_bF_buf86), .D(_3268_), .Q(micro_hash_synth_2_W_4__7_) );
	DFFPOSX1 DFFPOSX1_257 ( .CLK(clk_bF_buf85), .D(_3225_), .Q(micro_hash_synth_2_W_23__0_) );
	DFFPOSX1 DFFPOSX1_258 ( .CLK(clk_bF_buf84), .D(_3226_), .Q(micro_hash_synth_2_W_23__1_) );
	DFFPOSX1 DFFPOSX1_259 ( .CLK(clk_bF_buf83), .D(_3227_), .Q(micro_hash_synth_2_W_23__2_) );
	DFFPOSX1 DFFPOSX1_260 ( .CLK(clk_bF_buf82), .D(_3228_), .Q(micro_hash_synth_2_W_23__3_) );
	DFFPOSX1 DFFPOSX1_261 ( .CLK(clk_bF_buf81), .D(_3229_), .Q(micro_hash_synth_2_W_23__4_) );
	DFFPOSX1 DFFPOSX1_262 ( .CLK(clk_bF_buf80), .D(_3230_), .Q(micro_hash_synth_2_W_23__5_) );
	DFFPOSX1 DFFPOSX1_263 ( .CLK(clk_bF_buf79), .D(_3231_), .Q(micro_hash_synth_2_W_23__6_) );
	DFFPOSX1 DFFPOSX1_264 ( .CLK(clk_bF_buf78), .D(_3232_), .Q(micro_hash_synth_2_W_23__7_) );
	DFFPOSX1 DFFPOSX1_265 ( .CLK(clk_bF_buf77), .D(_3216_), .Q(micro_hash_synth_2_W_24__0_) );
	DFFPOSX1 DFFPOSX1_266 ( .CLK(clk_bF_buf76), .D(_3217_), .Q(micro_hash_synth_2_W_24__1_) );
	DFFPOSX1 DFFPOSX1_267 ( .CLK(clk_bF_buf75), .D(_3218_), .Q(micro_hash_synth_2_W_24__2_) );
	DFFPOSX1 DFFPOSX1_268 ( .CLK(clk_bF_buf74), .D(_3219_), .Q(micro_hash_synth_2_W_24__3_) );
	DFFPOSX1 DFFPOSX1_269 ( .CLK(clk_bF_buf73), .D(_3220_), .Q(micro_hash_synth_2_W_24__4_) );
	DFFPOSX1 DFFPOSX1_270 ( .CLK(clk_bF_buf72), .D(_3221_), .Q(micro_hash_synth_2_W_24__5_) );
	DFFPOSX1 DFFPOSX1_271 ( .CLK(clk_bF_buf71), .D(_3223_), .Q(micro_hash_synth_2_W_24__6_) );
	DFFPOSX1 DFFPOSX1_272 ( .CLK(clk_bF_buf70), .D(_3224_), .Q(micro_hash_synth_2_W_24__7_) );
	DFFPOSX1 DFFPOSX1_273 ( .CLK(clk_bF_buf69), .D(_3244_), .Q(micro_hash_synth_2_W_25__0_) );
	DFFPOSX1 DFFPOSX1_274 ( .CLK(clk_bF_buf68), .D(_3255_), .Q(micro_hash_synth_2_W_25__1_) );
	DFFPOSX1 DFFPOSX1_275 ( .CLK(clk_bF_buf67), .D(_3266_), .Q(micro_hash_synth_2_W_25__2_) );
	DFFPOSX1 DFFPOSX1_276 ( .CLK(clk_bF_buf66), .D(_3277_), .Q(micro_hash_synth_2_W_25__3_) );
	DFFPOSX1 DFFPOSX1_277 ( .CLK(clk_bF_buf65), .D(_3288_), .Q(micro_hash_synth_2_W_25__4_) );
	DFFPOSX1 DFFPOSX1_278 ( .CLK(clk_bF_buf64), .D(_3295_), .Q(micro_hash_synth_2_W_25__5_) );
	DFFPOSX1 DFFPOSX1_279 ( .CLK(clk_bF_buf63), .D(_3296_), .Q(micro_hash_synth_2_W_25__6_) );
	DFFPOSX1 DFFPOSX1_280 ( .CLK(clk_bF_buf62), .D(_3297_), .Q(micro_hash_synth_2_W_25__7_) );
	DFFPOSX1 DFFPOSX1_281 ( .CLK(clk_bF_buf61), .D(_3210_), .Q(micro_hash_synth_2_W_26__0_) );
	DFFPOSX1 DFFPOSX1_282 ( .CLK(clk_bF_buf60), .D(_3211_), .Q(micro_hash_synth_2_W_26__1_) );
	DFFPOSX1 DFFPOSX1_283 ( .CLK(clk_bF_buf59), .D(_3212_), .Q(micro_hash_synth_2_W_26__2_) );
	DFFPOSX1 DFFPOSX1_284 ( .CLK(clk_bF_buf58), .D(_3213_), .Q(micro_hash_synth_2_W_26__3_) );
	DFFPOSX1 DFFPOSX1_285 ( .CLK(clk_bF_buf57), .D(_3214_), .Q(micro_hash_synth_2_W_26__4_) );
	DFFPOSX1 DFFPOSX1_286 ( .CLK(clk_bF_buf56), .D(_3215_), .Q(micro_hash_synth_2_W_26__5_) );
	DFFPOSX1 DFFPOSX1_287 ( .CLK(clk_bF_buf55), .D(_3222_), .Q(micro_hash_synth_2_W_26__6_) );
	DFFPOSX1 DFFPOSX1_288 ( .CLK(clk_bF_buf54), .D(_3233_), .Q(micro_hash_synth_2_W_26__7_) );
	DFFPOSX1 DFFPOSX1_289 ( .CLK(clk_bF_buf53), .D(_3170_), .Q(micro_hash_synth_2_W_27__0_) );
	DFFPOSX1 DFFPOSX1_290 ( .CLK(clk_bF_buf52), .D(_3171_), .Q(micro_hash_synth_2_W_27__1_) );
	DFFPOSX1 DFFPOSX1_291 ( .CLK(clk_bF_buf51), .D(_3172_), .Q(micro_hash_synth_2_W_27__2_) );
	DFFPOSX1 DFFPOSX1_292 ( .CLK(clk_bF_buf50), .D(_3173_), .Q(micro_hash_synth_2_W_27__3_) );
	DFFPOSX1 DFFPOSX1_293 ( .CLK(clk_bF_buf49), .D(_3174_), .Q(micro_hash_synth_2_W_27__4_) );
	DFFPOSX1 DFFPOSX1_294 ( .CLK(clk_bF_buf48), .D(_3175_), .Q(micro_hash_synth_2_W_27__5_) );
	DFFPOSX1 DFFPOSX1_295 ( .CLK(clk_bF_buf47), .D(_3176_), .Q(micro_hash_synth_2_W_27__6_) );
	DFFPOSX1 DFFPOSX1_296 ( .CLK(clk_bF_buf46), .D(_3177_), .Q(micro_hash_synth_2_W_27__7_) );
	DFFPOSX1 DFFPOSX1_297 ( .CLK(clk_bF_buf45), .D(_3178_), .Q(micro_hash_synth_2_W_28__0_) );
	DFFPOSX1 DFFPOSX1_298 ( .CLK(clk_bF_buf44), .D(_3179_), .Q(micro_hash_synth_2_W_28__1_) );
	DFFPOSX1 DFFPOSX1_299 ( .CLK(clk_bF_buf43), .D(_3180_), .Q(micro_hash_synth_2_W_28__2_) );
	DFFPOSX1 DFFPOSX1_300 ( .CLK(clk_bF_buf42), .D(_3181_), .Q(micro_hash_synth_2_W_28__3_) );
	DFFPOSX1 DFFPOSX1_301 ( .CLK(clk_bF_buf41), .D(_3182_), .Q(micro_hash_synth_2_W_28__4_) );
	DFFPOSX1 DFFPOSX1_302 ( .CLK(clk_bF_buf40), .D(_3183_), .Q(micro_hash_synth_2_W_28__5_) );
	DFFPOSX1 DFFPOSX1_303 ( .CLK(clk_bF_buf39), .D(_3184_), .Q(micro_hash_synth_2_W_28__6_) );
	DFFPOSX1 DFFPOSX1_304 ( .CLK(clk_bF_buf38), .D(_3185_), .Q(micro_hash_synth_2_W_28__7_) );
	DFFPOSX1 DFFPOSX1_305 ( .CLK(clk_bF_buf37), .D(_3186_), .Q(micro_hash_synth_2_W_29__0_) );
	DFFPOSX1 DFFPOSX1_306 ( .CLK(clk_bF_buf36), .D(_3187_), .Q(micro_hash_synth_2_W_29__1_) );
	DFFPOSX1 DFFPOSX1_307 ( .CLK(clk_bF_buf35), .D(_3188_), .Q(micro_hash_synth_2_W_29__2_) );
	DFFPOSX1 DFFPOSX1_308 ( .CLK(clk_bF_buf34), .D(_3189_), .Q(micro_hash_synth_2_W_29__3_) );
	DFFPOSX1 DFFPOSX1_309 ( .CLK(clk_bF_buf33), .D(_3190_), .Q(micro_hash_synth_2_W_29__4_) );
	DFFPOSX1 DFFPOSX1_310 ( .CLK(clk_bF_buf32), .D(_3191_), .Q(micro_hash_synth_2_W_29__5_) );
	DFFPOSX1 DFFPOSX1_311 ( .CLK(clk_bF_buf31), .D(_3192_), .Q(micro_hash_synth_2_W_29__6_) );
	DFFPOSX1 DFFPOSX1_312 ( .CLK(clk_bF_buf30), .D(_3193_), .Q(micro_hash_synth_2_W_29__7_) );
	DFFPOSX1 DFFPOSX1_313 ( .CLK(clk_bF_buf29), .D(_3194_), .Q(micro_hash_synth_2_W_30__0_) );
	DFFPOSX1 DFFPOSX1_314 ( .CLK(clk_bF_buf28), .D(_3195_), .Q(micro_hash_synth_2_W_30__1_) );
	DFFPOSX1 DFFPOSX1_315 ( .CLK(clk_bF_buf27), .D(_3196_), .Q(micro_hash_synth_2_W_30__2_) );
	DFFPOSX1 DFFPOSX1_316 ( .CLK(clk_bF_buf26), .D(_3197_), .Q(micro_hash_synth_2_W_30__3_) );
	DFFPOSX1 DFFPOSX1_317 ( .CLK(clk_bF_buf25), .D(_3198_), .Q(micro_hash_synth_2_W_30__4_) );
	DFFPOSX1 DFFPOSX1_318 ( .CLK(clk_bF_buf24), .D(_3199_), .Q(micro_hash_synth_2_W_30__5_) );
	DFFPOSX1 DFFPOSX1_319 ( .CLK(clk_bF_buf23), .D(_3200_), .Q(micro_hash_synth_2_W_30__6_) );
	DFFPOSX1 DFFPOSX1_320 ( .CLK(clk_bF_buf22), .D(_3201_), .Q(micro_hash_synth_2_W_30__7_) );
	DFFPOSX1 DFFPOSX1_321 ( .CLK(clk_bF_buf21), .D(_3066_), .Q(micro_hash_synth_2_W_3__0_) );
	DFFPOSX1 DFFPOSX1_322 ( .CLK(clk_bF_buf20), .D(_3067_), .Q(micro_hash_synth_2_W_3__1_) );
	DFFPOSX1 DFFPOSX1_323 ( .CLK(clk_bF_buf19), .D(_3076_), .Q(micro_hash_synth_2_W_3__2_) );
	DFFPOSX1 DFFPOSX1_324 ( .CLK(clk_bF_buf18), .D(_3079_), .Q(micro_hash_synth_2_W_3__3_) );
	DFFPOSX1 DFFPOSX1_325 ( .CLK(clk_bF_buf17), .D(_3095_), .Q(micro_hash_synth_2_W_3__4_) );
	DFFPOSX1 DFFPOSX1_326 ( .CLK(clk_bF_buf16), .D(_3111_), .Q(micro_hash_synth_2_W_3__5_) );
	DFFPOSX1 DFFPOSX1_327 ( .CLK(clk_bF_buf15), .D(_3127_), .Q(micro_hash_synth_2_W_3__6_) );
	DFFPOSX1 DFFPOSX1_328 ( .CLK(clk_bF_buf14), .D(_3143_), .Q(micro_hash_synth_2_W_3__7_) );
	DFFPOSX1 DFFPOSX1_329 ( .CLK(clk_bF_buf13), .D(_3202_), .Q(micro_hash_synth_2_W_31__0_) );
	DFFPOSX1 DFFPOSX1_330 ( .CLK(clk_bF_buf12), .D(_3203_), .Q(micro_hash_synth_2_W_31__1_) );
	DFFPOSX1 DFFPOSX1_331 ( .CLK(clk_bF_buf11), .D(_3204_), .Q(micro_hash_synth_2_W_31__2_) );
	DFFPOSX1 DFFPOSX1_332 ( .CLK(clk_bF_buf10), .D(_3205_), .Q(micro_hash_synth_2_W_31__3_) );
	DFFPOSX1 DFFPOSX1_333 ( .CLK(clk_bF_buf9), .D(_3206_), .Q(micro_hash_synth_2_W_31__4_) );
	DFFPOSX1 DFFPOSX1_334 ( .CLK(clk_bF_buf8), .D(_3207_), .Q(micro_hash_synth_2_W_31__5_) );
	DFFPOSX1 DFFPOSX1_335 ( .CLK(clk_bF_buf7), .D(_3208_), .Q(micro_hash_synth_2_W_31__6_) );
	DFFPOSX1 DFFPOSX1_336 ( .CLK(clk_bF_buf6), .D(_3209_), .Q(micro_hash_synth_2_W_31__7_) );
	DFFPOSX1 DFFPOSX1_337 ( .CLK(clk_bF_buf5), .D(_3137_), .Q(micro_hash_synth_2_W_1__0_) );
	DFFPOSX1 DFFPOSX1_338 ( .CLK(clk_bF_buf4), .D(_3138_), .Q(micro_hash_synth_2_W_1__1_) );
	DFFPOSX1 DFFPOSX1_339 ( .CLK(clk_bF_buf3), .D(_3139_), .Q(micro_hash_synth_2_W_1__2_) );
	DFFPOSX1 DFFPOSX1_340 ( .CLK(clk_bF_buf2), .D(_3140_), .Q(micro_hash_synth_2_W_1__3_) );
	DFFPOSX1 DFFPOSX1_341 ( .CLK(clk_bF_buf1), .D(_3141_), .Q(micro_hash_synth_2_W_1__4_) );
	DFFPOSX1 DFFPOSX1_342 ( .CLK(clk_bF_buf0), .D(_3142_), .Q(micro_hash_synth_2_W_1__5_) );
	DFFPOSX1 DFFPOSX1_343 ( .CLK(clk_bF_buf113), .D(_3144_), .Q(micro_hash_synth_2_W_1__6_) );
	DFFPOSX1 DFFPOSX1_344 ( .CLK(clk_bF_buf112), .D(_3145_), .Q(micro_hash_synth_2_W_1__7_) );
	DFFPOSX1 DFFPOSX1_345 ( .CLK(clk_bF_buf111), .D(_3162_), .Q(micro_hash_synth_2_W_2__0_) );
	DFFPOSX1 DFFPOSX1_346 ( .CLK(clk_bF_buf110), .D(_3163_), .Q(micro_hash_synth_2_W_2__1_) );
	DFFPOSX1 DFFPOSX1_347 ( .CLK(clk_bF_buf109), .D(_3164_), .Q(micro_hash_synth_2_W_2__2_) );
	DFFPOSX1 DFFPOSX1_348 ( .CLK(clk_bF_buf108), .D(_3165_), .Q(micro_hash_synth_2_W_2__3_) );
	DFFPOSX1 DFFPOSX1_349 ( .CLK(clk_bF_buf107), .D(_3166_), .Q(micro_hash_synth_2_W_2__4_) );
	DFFPOSX1 DFFPOSX1_350 ( .CLK(clk_bF_buf106), .D(_3167_), .Q(micro_hash_synth_2_W_2__5_) );
	DFFPOSX1 DFFPOSX1_351 ( .CLK(clk_bF_buf105), .D(_3168_), .Q(micro_hash_synth_2_W_2__6_) );
	DFFPOSX1 DFFPOSX1_352 ( .CLK(clk_bF_buf104), .D(_3169_), .Q(micro_hash_synth_2_W_2__7_) );
	NOR2X1 NOR2X1_94 ( .A(concatenador_counter_2_), .B(concatenador_counter_1_bF_buf7), .Y(_4906_) );
	NAND2X1 NAND2X1_190 ( .A(concatenador_counter_5_), .B(concatenador_counter_0_bF_buf13), .Y(_4907_) );
	NOR3X1 NOR3X1_1 ( .A(concatenador_counter_4_), .B(concatenador_counter_3_), .C(_4907_), .Y(_4908_) );
	AOI21X1 AOI21X1_175 ( .A(_4906_), .B(_4908_), .C(mux0_sel_bF_buf5), .Y(_4909_) );
	OR2X2 OR2X2_11 ( .A(concatenador_counter_2d_2_), .B(concatenador_counter_2d_1_bF_buf2), .Y(_4910_) );
	OR2X2 OR2X2_12 ( .A(concatenador_counter_2d_4_), .B(concatenador_counter_2d_3_), .Y(_4911_) );
	NAND2X1 NAND2X1_191 ( .A(concatenador_counter_2d_5_), .B(concatenador_counter_2d_0_bF_buf10), .Y(_4912_) );
	NOR3X1 NOR3X1_2 ( .A(_4910_), .B(_4912_), .C(_4911_), .Y(_4913_) );
	OAI21X1 OAI21X1_333 ( .A(_4909_), .B(_4913_), .C(reset_L_bF_buf48), .Y(_4858_) );
	INVX1 INVX1_272 ( .A(Hhash_synth2_0_), .Y(_4914_) );
	INVX2 INVX2_2 ( .A(reset_L_bF_buf47), .Y(_4915_) );
	AOI21X1 AOI21X1_176 ( .A(mux0_sel_bF_buf4), .B(Hhash_synth1_0_), .C(_4915_), .Y(_4916_) );
	OAI21X1 OAI21X1_334 ( .A(mux0_sel_bF_buf3), .B(_4914_), .C(_4916_), .Y(_4857__0_) );
	NOR2X1 NOR2X1_95 ( .A(mux0_sel_bF_buf2), .B(Hhash_synth2_1_), .Y(_4859_) );
	INVX4 INVX4_1 ( .A(mux0_sel_bF_buf1), .Y(_4860_) );
	OAI21X1 OAI21X1_335 ( .A(_4860_), .B(Hhash_synth1_1_), .C(reset_L_bF_buf46), .Y(_4861_) );
	NOR2X1 NOR2X1_96 ( .A(_4859_), .B(_4861_), .Y(_4857__1_) );
	NOR2X1 NOR2X1_97 ( .A(mux0_sel_bF_buf0), .B(Hhash_synth2_2_), .Y(_4862_) );
	OAI21X1 OAI21X1_336 ( .A(_4860_), .B(Hhash_synth1_2_), .C(reset_L_bF_buf45), .Y(_4863_) );
	NOR2X1 NOR2X1_98 ( .A(_4862_), .B(_4863_), .Y(_4857__2_) );
	NOR2X1 NOR2X1_99 ( .A(mux0_sel_bF_buf5), .B(Hhash_synth2_3_), .Y(_4864_) );
	OAI21X1 OAI21X1_337 ( .A(_4860_), .B(Hhash_synth1_3_), .C(reset_L_bF_buf44), .Y(_4865_) );
	NOR2X1 NOR2X1_100 ( .A(_4864_), .B(_4865_), .Y(_4857__3_) );
	NOR2X1 NOR2X1_101 ( .A(mux0_sel_bF_buf4), .B(Hhash_synth2_4_), .Y(_4866_) );
	OAI21X1 OAI21X1_338 ( .A(_4860_), .B(Hhash_synth1_4_), .C(reset_L_bF_buf43), .Y(_4867_) );
	NOR2X1 NOR2X1_102 ( .A(_4866_), .B(_4867_), .Y(_4857__4_) );
	NOR2X1 NOR2X1_103 ( .A(mux0_sel_bF_buf3), .B(Hhash_synth2_5_), .Y(_4868_) );
	OAI21X1 OAI21X1_339 ( .A(_4860_), .B(Hhash_synth1_5_), .C(reset_L_bF_buf42), .Y(_4869_) );
	NOR2X1 NOR2X1_104 ( .A(_4868_), .B(_4869_), .Y(_4857__5_) );
	NOR2X1 NOR2X1_105 ( .A(mux0_sel_bF_buf2), .B(Hhash_synth2_6_), .Y(_4870_) );
	OAI21X1 OAI21X1_340 ( .A(_4860_), .B(Hhash_synth1_6_), .C(reset_L_bF_buf41), .Y(_4871_) );
	NOR2X1 NOR2X1_106 ( .A(_4870_), .B(_4871_), .Y(_4857__6_) );
	NOR2X1 NOR2X1_107 ( .A(mux0_sel_bF_buf1), .B(Hhash_synth2_7_), .Y(_4872_) );
	OAI21X1 OAI21X1_341 ( .A(_4860_), .B(Hhash_synth1_7_), .C(reset_L_bF_buf40), .Y(_4873_) );
	NOR2X1 NOR2X1_108 ( .A(_4872_), .B(_4873_), .Y(_4857__7_) );
	INVX1 INVX1_273 ( .A(Hhash_synth2_8_), .Y(_4874_) );
	AOI21X1 AOI21X1_177 ( .A(mux0_sel_bF_buf0), .B(Hhash_synth1_8_), .C(_4915_), .Y(_4875_) );
	OAI21X1 OAI21X1_342 ( .A(mux0_sel_bF_buf5), .B(_4874_), .C(_4875_), .Y(_4857__8_) );
	NOR2X1 NOR2X1_109 ( .A(mux0_sel_bF_buf4), .B(Hhash_synth2_9_), .Y(_4876_) );
	OAI21X1 OAI21X1_343 ( .A(_4860_), .B(Hhash_synth1_9_), .C(reset_L_bF_buf39), .Y(_4877_) );
	NOR2X1 NOR2X1_110 ( .A(_4876_), .B(_4877_), .Y(_4857__9_) );
	NOR2X1 NOR2X1_111 ( .A(mux0_sel_bF_buf3), .B(Hhash_synth2_10_), .Y(_4878_) );
	OAI21X1 OAI21X1_344 ( .A(_4860_), .B(Hhash_synth1_10_), .C(reset_L_bF_buf38), .Y(_4879_) );
	NOR2X1 NOR2X1_112 ( .A(_4878_), .B(_4879_), .Y(_4857__10_) );
	INVX1 INVX1_274 ( .A(Hhash_synth2_11_), .Y(_4880_) );
	AOI21X1 AOI21X1_178 ( .A(mux0_sel_bF_buf2), .B(Hhash_synth1_11_), .C(_4915_), .Y(_4881_) );
	OAI21X1 OAI21X1_345 ( .A(mux0_sel_bF_buf1), .B(_4880_), .C(_4881_), .Y(_4857__11_) );
	NOR2X1 NOR2X1_113 ( .A(mux0_sel_bF_buf0), .B(Hhash_synth2_12_), .Y(_4882_) );
	OAI21X1 OAI21X1_346 ( .A(_4860_), .B(Hhash_synth1_12_), .C(reset_L_bF_buf37), .Y(_4883_) );
	NOR2X1 NOR2X1_114 ( .A(_4882_), .B(_4883_), .Y(_4857__12_) );
	NOR2X1 NOR2X1_115 ( .A(mux0_sel_bF_buf5), .B(Hhash_synth2_13_), .Y(_4884_) );
	OAI21X1 OAI21X1_347 ( .A(_4860_), .B(Hhash_synth1_13_), .C(reset_L_bF_buf36), .Y(_4885_) );
	NOR2X1 NOR2X1_116 ( .A(_4884_), .B(_4885_), .Y(_4857__13_) );
	NOR2X1 NOR2X1_117 ( .A(mux0_sel_bF_buf4), .B(Hhash_synth2_14_), .Y(_4886_) );
	OAI21X1 OAI21X1_348 ( .A(_4860_), .B(Hhash_synth1_14_), .C(reset_L_bF_buf35), .Y(_4887_) );
	NOR2X1 NOR2X1_118 ( .A(_4886_), .B(_4887_), .Y(_4857__14_) );
	INVX1 INVX1_275 ( .A(Hhash_synth2_15_), .Y(_4888_) );
	AOI21X1 AOI21X1_179 ( .A(mux0_sel_bF_buf3), .B(Hhash_synth1_15_), .C(_4915_), .Y(_4889_) );
	OAI21X1 OAI21X1_349 ( .A(mux0_sel_bF_buf2), .B(_4888_), .C(_4889_), .Y(_4857__15_) );
	NOR2X1 NOR2X1_119 ( .A(mux0_sel_bF_buf1), .B(Hhash_synth2_16_), .Y(_4890_) );
	OAI21X1 OAI21X1_350 ( .A(_4860_), .B(Hhash_synth1_16_), .C(reset_L_bF_buf34), .Y(_4891_) );
	NOR2X1 NOR2X1_120 ( .A(_4890_), .B(_4891_), .Y(_4857__16_) );
	INVX1 INVX1_276 ( .A(Hhash_synth2_17_), .Y(_4892_) );
	AOI21X1 AOI21X1_180 ( .A(mux0_sel_bF_buf0), .B(Hhash_synth1_17_), .C(_4915_), .Y(_4893_) );
	OAI21X1 OAI21X1_351 ( .A(mux0_sel_bF_buf5), .B(_4892_), .C(_4893_), .Y(_4857__17_) );
	INVX1 INVX1_277 ( .A(Hhash_synth2_18_), .Y(_4894_) );
	AOI21X1 AOI21X1_181 ( .A(mux0_sel_bF_buf4), .B(Hhash_synth1_18_), .C(_4915_), .Y(_4895_) );
	OAI21X1 OAI21X1_352 ( .A(mux0_sel_bF_buf3), .B(_4894_), .C(_4895_), .Y(_4857__18_) );
	INVX1 INVX1_278 ( .A(Hhash_synth2_19_), .Y(_4896_) );
	AOI21X1 AOI21X1_182 ( .A(mux0_sel_bF_buf2), .B(Hhash_synth1_19_), .C(_4915_), .Y(_4897_) );
	OAI21X1 OAI21X1_353 ( .A(mux0_sel_bF_buf1), .B(_4896_), .C(_4897_), .Y(_4857__19_) );
	INVX1 INVX1_279 ( .A(Hhash_synth2_20_), .Y(_4898_) );
	AOI21X1 AOI21X1_183 ( .A(mux0_sel_bF_buf0), .B(Hhash_synth1_20_), .C(_4915_), .Y(_4899_) );
	OAI21X1 OAI21X1_354 ( .A(mux0_sel_bF_buf5), .B(_4898_), .C(_4899_), .Y(_4857__20_) );
	INVX1 INVX1_280 ( .A(Hhash_synth2_21_), .Y(_4900_) );
	AOI21X1 AOI21X1_184 ( .A(mux0_sel_bF_buf4), .B(Hhash_synth1_21_), .C(_4915_), .Y(_4901_) );
	OAI21X1 OAI21X1_355 ( .A(mux0_sel_bF_buf3), .B(_4900_), .C(_4901_), .Y(_4857__21_) );
	INVX1 INVX1_281 ( .A(Hhash_synth2_22_), .Y(_4902_) );
	AOI21X1 AOI21X1_185 ( .A(mux0_sel_bF_buf2), .B(Hhash_synth1_22_), .C(_4915_), .Y(_4903_) );
	OAI21X1 OAI21X1_356 ( .A(mux0_sel_bF_buf1), .B(_4902_), .C(_4903_), .Y(_4857__22_) );
	INVX1 INVX1_282 ( .A(Hhash_synth2_23_), .Y(_4904_) );
	AOI21X1 AOI21X1_186 ( .A(mux0_sel_bF_buf0), .B(Hhash_synth1_23_), .C(_4915_), .Y(_4905_) );
	OAI21X1 OAI21X1_357 ( .A(mux0_sel_bF_buf5), .B(_4904_), .C(_4905_), .Y(_4857__23_) );
	DFFPOSX1 DFFPOSX1_353 ( .CLK(clk_bF_buf103), .D(_4857__0_), .Q(Y_0_) );
	DFFPOSX1 DFFPOSX1_354 ( .CLK(clk_bF_buf102), .D(_4857__1_), .Q(Y_1_) );
	DFFPOSX1 DFFPOSX1_355 ( .CLK(clk_bF_buf101), .D(_4857__2_), .Q(Y_2_) );
	DFFPOSX1 DFFPOSX1_356 ( .CLK(clk_bF_buf100), .D(_4857__3_), .Q(Y_3_) );
	DFFPOSX1 DFFPOSX1_357 ( .CLK(clk_bF_buf99), .D(_4857__4_), .Q(Y_4_) );
	DFFPOSX1 DFFPOSX1_358 ( .CLK(clk_bF_buf98), .D(_4857__5_), .Q(Y_5_) );
	DFFPOSX1 DFFPOSX1_359 ( .CLK(clk_bF_buf97), .D(_4857__6_), .Q(Y_6_) );
	DFFPOSX1 DFFPOSX1_360 ( .CLK(clk_bF_buf96), .D(_4857__7_), .Q(Y_7_) );
	DFFPOSX1 DFFPOSX1_361 ( .CLK(clk_bF_buf95), .D(_4857__8_), .Q(Y_8_) );
	DFFPOSX1 DFFPOSX1_362 ( .CLK(clk_bF_buf94), .D(_4857__9_), .Q(Y_9_) );
	DFFPOSX1 DFFPOSX1_363 ( .CLK(clk_bF_buf93), .D(_4857__10_), .Q(Y_10_) );
	DFFPOSX1 DFFPOSX1_364 ( .CLK(clk_bF_buf92), .D(_4857__11_), .Q(Y_11_) );
	DFFPOSX1 DFFPOSX1_365 ( .CLK(clk_bF_buf91), .D(_4857__12_), .Q(Y_12_) );
	DFFPOSX1 DFFPOSX1_366 ( .CLK(clk_bF_buf90), .D(_4857__13_), .Q(Y_13_) );
	DFFPOSX1 DFFPOSX1_367 ( .CLK(clk_bF_buf89), .D(_4857__14_), .Q(Y_14_) );
	DFFPOSX1 DFFPOSX1_368 ( .CLK(clk_bF_buf88), .D(_4857__15_), .Q(Y_15_) );
	DFFPOSX1 DFFPOSX1_369 ( .CLK(clk_bF_buf87), .D(_4857__16_), .Q(Y_16_) );
	DFFPOSX1 DFFPOSX1_370 ( .CLK(clk_bF_buf86), .D(_4857__17_), .Q(Y_17_) );
	DFFPOSX1 DFFPOSX1_371 ( .CLK(clk_bF_buf85), .D(_4857__18_), .Q(Y_18_) );
	DFFPOSX1 DFFPOSX1_372 ( .CLK(clk_bF_buf84), .D(_4857__19_), .Q(Y_19_) );
	DFFPOSX1 DFFPOSX1_373 ( .CLK(clk_bF_buf83), .D(_4857__20_), .Q(Y_20_) );
	DFFPOSX1 DFFPOSX1_374 ( .CLK(clk_bF_buf82), .D(_4857__21_), .Q(Y_21_) );
	DFFPOSX1 DFFPOSX1_375 ( .CLK(clk_bF_buf81), .D(_4857__22_), .Q(Y_22_) );
	DFFPOSX1 DFFPOSX1_376 ( .CLK(clk_bF_buf80), .D(_4857__23_), .Q(Y_23_) );
	DFFPOSX1 DFFPOSX1_377 ( .CLK(clk_bF_buf79), .D(_4858_), .Q(mux0_sel) );
	INVX8 INVX8_2 ( .A(mux1_sel_bF_buf4), .Y(_4919_) );
	NOR2X1 NOR2X1_121 ( .A(concatenador_counter_1_bF_buf6), .B(concatenador_counter_0_bF_buf12), .Y(_4920_) );
	NOR2X1 NOR2X1_122 ( .A(concatenador_counter_3_), .B(concatenador_counter_2_), .Y(_4921_) );
	NOR2X1 NOR2X1_123 ( .A(concatenador_counter_5_), .B(concatenador_counter_4_), .Y(_4922_) );
	NAND3X1 NAND3X1_57 ( .A(_4920_), .B(_4921_), .C(_4922_), .Y(_4923_) );
	AND2X2 AND2X2_31 ( .A(_4923_), .B(_4919__bF_buf4), .Y(_4924_) );
	OR2X2 OR2X2_13 ( .A(concatenador_counter_2d_1_bF_buf1), .B(concatenador_counter_2d_0_bF_buf9), .Y(_4925_) );
	OR2X2 OR2X2_14 ( .A(concatenador_counter_2d_2_), .B(concatenador_counter_2d_5_), .Y(_4926_) );
	OR2X2 OR2X2_15 ( .A(concatenador_counter_2d_3_), .B(concatenador_counter_2d_4_), .Y(_4927_) );
	NOR3X1 NOR3X1_3 ( .A(_4925_), .B(_4926_), .C(_4927_), .Y(_4928_) );
	OAI21X1 OAI21X1_358 ( .A(_4924_), .B(_4928_), .C(reset_L_bF_buf33), .Y(_4918_) );
	NOR2X1 NOR2X1_124 ( .A(mux1_sel_bF_buf3), .B(micro_hash_synth_2_nonce_synth_1_0_), .Y(_4929_) );
	OAI21X1 OAI21X1_359 ( .A(_4919__bF_buf3), .B(micro_hash_synth_1_nonce_synth_1_0_), .C(reset_L_bF_buf32), .Y(_4930_) );
	NOR2X1 NOR2X1_125 ( .A(_4929_), .B(_4930_), .Y(_4917__0_) );
	NOR2X1 NOR2X1_126 ( .A(mux1_sel_bF_buf2), .B(micro_hash_synth_2_nonce_synth_1_1_), .Y(_4931_) );
	OAI21X1 OAI21X1_360 ( .A(_4919__bF_buf2), .B(micro_hash_synth_1_nonce_synth_1_1_), .C(reset_L_bF_buf31), .Y(_4932_) );
	NOR2X1 NOR2X1_127 ( .A(_4931_), .B(_4932_), .Y(_4917__1_) );
	NOR2X1 NOR2X1_128 ( .A(mux1_sel_bF_buf1), .B(micro_hash_synth_2_nonce_synth_1_2_), .Y(_4933_) );
	OAI21X1 OAI21X1_361 ( .A(_4919__bF_buf1), .B(micro_hash_synth_1_nonce_synth_1_2_), .C(reset_L_bF_buf30), .Y(_4934_) );
	NOR2X1 NOR2X1_129 ( .A(_4933_), .B(_4934_), .Y(_4917__2_) );
	NOR2X1 NOR2X1_130 ( .A(mux1_sel_bF_buf0), .B(micro_hash_synth_2_nonce_synth_1_3_), .Y(_4935_) );
	OAI21X1 OAI21X1_362 ( .A(_4919__bF_buf0), .B(micro_hash_synth_1_nonce_synth_1_3_), .C(reset_L_bF_buf29), .Y(_4936_) );
	NOR2X1 NOR2X1_131 ( .A(_4935_), .B(_4936_), .Y(_4917__3_) );
	NOR2X1 NOR2X1_132 ( .A(mux1_sel_bF_buf4), .B(micro_hash_synth_2_nonce_synth_1_4_), .Y(_4937_) );
	OAI21X1 OAI21X1_363 ( .A(_4919__bF_buf4), .B(micro_hash_synth_1_nonce_synth_1_4_), .C(reset_L_bF_buf28), .Y(_4938_) );
	NOR2X1 NOR2X1_133 ( .A(_4937_), .B(_4938_), .Y(_4917__4_) );
	NOR2X1 NOR2X1_134 ( .A(mux1_sel_bF_buf3), .B(micro_hash_synth_2_nonce_synth_1_5_), .Y(_4939_) );
	OAI21X1 OAI21X1_364 ( .A(_4919__bF_buf3), .B(micro_hash_synth_1_nonce_synth_1_5_), .C(reset_L_bF_buf27), .Y(_4940_) );
	NOR2X1 NOR2X1_135 ( .A(_4939_), .B(_4940_), .Y(_4917__5_) );
	NOR2X1 NOR2X1_136 ( .A(mux1_sel_bF_buf2), .B(micro_hash_synth_2_nonce_synth_1_6_), .Y(_4941_) );
	OAI21X1 OAI21X1_365 ( .A(_4919__bF_buf2), .B(micro_hash_synth_1_nonce_synth_1_6_), .C(reset_L_bF_buf26), .Y(_4942_) );
	NOR2X1 NOR2X1_137 ( .A(_4941_), .B(_4942_), .Y(_4917__6_) );
	NOR2X1 NOR2X1_138 ( .A(mux1_sel_bF_buf1), .B(micro_hash_synth_2_nonce_synth_1_7_), .Y(_4943_) );
	OAI21X1 OAI21X1_366 ( .A(_4919__bF_buf1), .B(micro_hash_synth_1_nonce_synth_1_7_), .C(reset_L_bF_buf25), .Y(_4944_) );
	NOR2X1 NOR2X1_139 ( .A(_4943_), .B(_4944_), .Y(_4917__7_) );
	NOR2X1 NOR2X1_140 ( .A(mux1_sel_bF_buf0), .B(micro_hash_synth_2_nonce_synth_1_8_), .Y(_4945_) );
	OAI21X1 OAI21X1_367 ( .A(_4919__bF_buf0), .B(micro_hash_synth_1_nonce_synth_1_8_), .C(reset_L_bF_buf24), .Y(_4946_) );
	NOR2X1 NOR2X1_141 ( .A(_4945_), .B(_4946_), .Y(_4917__8_) );
	NOR2X1 NOR2X1_142 ( .A(mux1_sel_bF_buf4), .B(micro_hash_synth_2_nonce_synth_1_9_), .Y(_4947_) );
	OAI21X1 OAI21X1_368 ( .A(_4919__bF_buf4), .B(micro_hash_synth_1_nonce_synth_1_9_), .C(reset_L_bF_buf23), .Y(_4948_) );
	NOR2X1 NOR2X1_143 ( .A(_4947_), .B(_4948_), .Y(_4917__9_) );
	NOR2X1 NOR2X1_144 ( .A(mux1_sel_bF_buf3), .B(micro_hash_synth_2_nonce_synth_1_10_), .Y(_4949_) );
	OAI21X1 OAI21X1_369 ( .A(_4919__bF_buf3), .B(micro_hash_synth_1_nonce_synth_1_10_), .C(reset_L_bF_buf22), .Y(_4950_) );
	NOR2X1 NOR2X1_145 ( .A(_4949_), .B(_4950_), .Y(_4917__10_) );
	NOR2X1 NOR2X1_146 ( .A(mux1_sel_bF_buf2), .B(micro_hash_synth_2_nonce_synth_1_11_), .Y(_4951_) );
	OAI21X1 OAI21X1_370 ( .A(_4919__bF_buf2), .B(micro_hash_synth_1_nonce_synth_1_11_), .C(reset_L_bF_buf21), .Y(_4952_) );
	NOR2X1 NOR2X1_147 ( .A(_4951_), .B(_4952_), .Y(_4917__11_) );
	NOR2X1 NOR2X1_148 ( .A(mux1_sel_bF_buf1), .B(micro_hash_synth_2_nonce_synth_1_12_), .Y(_4953_) );
	OAI21X1 OAI21X1_371 ( .A(_4919__bF_buf1), .B(micro_hash_synth_1_nonce_synth_1_12_), .C(reset_L_bF_buf20), .Y(_4954_) );
	NOR2X1 NOR2X1_149 ( .A(_4953_), .B(_4954_), .Y(_4917__12_) );
	NOR2X1 NOR2X1_150 ( .A(mux1_sel_bF_buf0), .B(micro_hash_synth_2_nonce_synth_1_13_), .Y(_4955_) );
	OAI21X1 OAI21X1_372 ( .A(_4919__bF_buf0), .B(micro_hash_synth_1_nonce_synth_1_13_), .C(reset_L_bF_buf19), .Y(_4956_) );
	NOR2X1 NOR2X1_151 ( .A(_4955_), .B(_4956_), .Y(_4917__13_) );
	NOR2X1 NOR2X1_152 ( .A(mux1_sel_bF_buf4), .B(micro_hash_synth_2_nonce_synth_1_14_), .Y(_4957_) );
	OAI21X1 OAI21X1_373 ( .A(_4919__bF_buf4), .B(micro_hash_synth_1_nonce_synth_1_14_), .C(reset_L_bF_buf18), .Y(_4958_) );
	NOR2X1 NOR2X1_153 ( .A(_4957_), .B(_4958_), .Y(_4917__14_) );
	NOR2X1 NOR2X1_154 ( .A(mux1_sel_bF_buf3), .B(micro_hash_synth_2_nonce_synth_1_15_), .Y(_4959_) );
	OAI21X1 OAI21X1_374 ( .A(_4919__bF_buf3), .B(micro_hash_synth_1_nonce_synth_1_15_), .C(reset_L_bF_buf17), .Y(_4960_) );
	NOR2X1 NOR2X1_155 ( .A(_4959_), .B(_4960_), .Y(_4917__15_) );
	NOR2X1 NOR2X1_156 ( .A(mux1_sel_bF_buf2), .B(micro_hash_synth_2_nonce_synth_1_16_), .Y(_4961_) );
	OAI21X1 OAI21X1_375 ( .A(_4919__bF_buf2), .B(micro_hash_synth_1_nonce_synth_1_16_), .C(reset_L_bF_buf16), .Y(_4962_) );
	NOR2X1 NOR2X1_157 ( .A(_4961_), .B(_4962_), .Y(_4917__16_) );
	NOR2X1 NOR2X1_158 ( .A(mux1_sel_bF_buf1), .B(micro_hash_synth_2_nonce_synth_1_17_), .Y(_4963_) );
	OAI21X1 OAI21X1_376 ( .A(_4919__bF_buf1), .B(micro_hash_synth_1_nonce_synth_1_17_), .C(reset_L_bF_buf15), .Y(_4964_) );
	NOR2X1 NOR2X1_159 ( .A(_4963_), .B(_4964_), .Y(_4917__17_) );
	NOR2X1 NOR2X1_160 ( .A(mux1_sel_bF_buf0), .B(micro_hash_synth_2_nonce_synth_1_18_), .Y(_4965_) );
	OAI21X1 OAI21X1_377 ( .A(_4919__bF_buf0), .B(micro_hash_synth_1_nonce_synth_1_18_), .C(reset_L_bF_buf14), .Y(_4966_) );
	NOR2X1 NOR2X1_161 ( .A(_4965_), .B(_4966_), .Y(_4917__18_) );
	NOR2X1 NOR2X1_162 ( .A(mux1_sel_bF_buf4), .B(micro_hash_synth_2_nonce_synth_1_19_), .Y(_4967_) );
	OAI21X1 OAI21X1_378 ( .A(_4919__bF_buf4), .B(micro_hash_synth_1_nonce_synth_1_19_), .C(reset_L_bF_buf13), .Y(_4968_) );
	NOR2X1 NOR2X1_163 ( .A(_4967_), .B(_4968_), .Y(_4917__19_) );
	NOR2X1 NOR2X1_164 ( .A(mux1_sel_bF_buf3), .B(micro_hash_synth_2_nonce_synth_1_20_), .Y(_4969_) );
	OAI21X1 OAI21X1_379 ( .A(_4919__bF_buf3), .B(micro_hash_synth_1_nonce_synth_1_20_), .C(reset_L_bF_buf12), .Y(_4970_) );
	NOR2X1 NOR2X1_165 ( .A(_4969_), .B(_4970_), .Y(_4917__20_) );
	NOR2X1 NOR2X1_166 ( .A(mux1_sel_bF_buf2), .B(micro_hash_synth_2_nonce_synth_1_21_), .Y(_4971_) );
	OAI21X1 OAI21X1_380 ( .A(_4919__bF_buf2), .B(micro_hash_synth_1_nonce_synth_1_21_), .C(reset_L_bF_buf11), .Y(_4972_) );
	NOR2X1 NOR2X1_167 ( .A(_4971_), .B(_4972_), .Y(_4917__21_) );
	NOR2X1 NOR2X1_168 ( .A(mux1_sel_bF_buf1), .B(micro_hash_synth_2_nonce_synth_1_22_), .Y(_4973_) );
	OAI21X1 OAI21X1_381 ( .A(_4919__bF_buf1), .B(micro_hash_synth_1_nonce_synth_1_22_), .C(reset_L_bF_buf10), .Y(_4974_) );
	NOR2X1 NOR2X1_169 ( .A(_4973_), .B(_4974_), .Y(_4917__22_) );
	NOR2X1 NOR2X1_170 ( .A(mux1_sel_bF_buf0), .B(micro_hash_synth_2_nonce_synth_1_23_), .Y(_4975_) );
	OAI21X1 OAI21X1_382 ( .A(_4919__bF_buf0), .B(micro_hash_synth_1_nonce_synth_1_23_), .C(reset_L_bF_buf9), .Y(_4976_) );
	NOR2X1 NOR2X1_171 ( .A(_4975_), .B(_4976_), .Y(_4917__23_) );
	NOR2X1 NOR2X1_172 ( .A(mux1_sel_bF_buf4), .B(micro_hash_synth_2_nonce_synth_1_24_), .Y(_4977_) );
	OAI21X1 OAI21X1_383 ( .A(_4919__bF_buf4), .B(micro_hash_synth_1_nonce_synth_1_24_), .C(reset_L_bF_buf8), .Y(_4978_) );
	NOR2X1 NOR2X1_173 ( .A(_4977_), .B(_4978_), .Y(_4917__24_) );
	NOR2X1 NOR2X1_174 ( .A(mux1_sel_bF_buf3), .B(micro_hash_synth_2_nonce_synth_1_25_), .Y(_4979_) );
	OAI21X1 OAI21X1_384 ( .A(_4919__bF_buf3), .B(micro_hash_synth_1_nonce_synth_1_25_), .C(reset_L_bF_buf7), .Y(_4980_) );
	NOR2X1 NOR2X1_175 ( .A(_4979_), .B(_4980_), .Y(_4917__25_) );
	NOR2X1 NOR2X1_176 ( .A(mux1_sel_bF_buf2), .B(micro_hash_synth_2_nonce_synth_1_26_), .Y(_4981_) );
	OAI21X1 OAI21X1_385 ( .A(_4919__bF_buf2), .B(micro_hash_synth_1_nonce_synth_1_26_), .C(reset_L_bF_buf6), .Y(_4982_) );
	NOR2X1 NOR2X1_177 ( .A(_4981_), .B(_4982_), .Y(_4917__26_) );
	NOR2X1 NOR2X1_178 ( .A(mux1_sel_bF_buf1), .B(micro_hash_synth_2_nonce_synth_1_27_), .Y(_4983_) );
	OAI21X1 OAI21X1_386 ( .A(_4919__bF_buf1), .B(micro_hash_synth_1_nonce_synth_1_27_), .C(reset_L_bF_buf5), .Y(_4984_) );
	NOR2X1 NOR2X1_179 ( .A(_4983_), .B(_4984_), .Y(_4917__27_) );
	NOR2X1 NOR2X1_180 ( .A(mux1_sel_bF_buf0), .B(micro_hash_synth_2_nonce_synth_1_28_), .Y(_4985_) );
	OAI21X1 OAI21X1_387 ( .A(_4919__bF_buf0), .B(micro_hash_synth_1_nonce_synth_1_28_), .C(reset_L_bF_buf4), .Y(_4986_) );
	NOR2X1 NOR2X1_181 ( .A(_4985_), .B(_4986_), .Y(_4917__28_) );
	NOR2X1 NOR2X1_182 ( .A(mux1_sel_bF_buf4), .B(micro_hash_synth_2_nonce_synth_1_29_), .Y(_4987_) );
	OAI21X1 OAI21X1_388 ( .A(_4919__bF_buf4), .B(micro_hash_synth_1_nonce_synth_1_29_), .C(reset_L_bF_buf3), .Y(_4988_) );
	NOR2X1 NOR2X1_183 ( .A(_4987_), .B(_4988_), .Y(_4917__29_) );
	NOR2X1 NOR2X1_184 ( .A(mux1_sel_bF_buf3), .B(micro_hash_synth_2_nonce_synth_1_30_), .Y(_4989_) );
	OAI21X1 OAI21X1_389 ( .A(_4919__bF_buf3), .B(micro_hash_synth_1_nonce_synth_1_30_), .C(reset_L_bF_buf2), .Y(_4990_) );
	NOR2X1 NOR2X1_185 ( .A(_4989_), .B(_4990_), .Y(_4917__30_) );
	NOR2X1 NOR2X1_186 ( .A(mux1_sel_bF_buf2), .B(micro_hash_synth_2_nonce_synth_1_31_), .Y(_4991_) );
	OAI21X1 OAI21X1_390 ( .A(_4919__bF_buf2), .B(micro_hash_synth_1_nonce_synth_1_31_), .C(reset_L_bF_buf1), .Y(_4992_) );
	NOR2X1 NOR2X1_187 ( .A(_4991_), .B(_4992_), .Y(_4917__31_) );
	DFFPOSX1 DFFPOSX1_378 ( .CLK(clk_bF_buf78), .D(_4917__0_), .Q(Ynonce_synth_0_) );
	DFFPOSX1 DFFPOSX1_379 ( .CLK(clk_bF_buf77), .D(_4917__1_), .Q(Ynonce_synth_1_) );
	DFFPOSX1 DFFPOSX1_380 ( .CLK(clk_bF_buf76), .D(_4917__2_), .Q(Ynonce_synth_2_) );
	DFFPOSX1 DFFPOSX1_381 ( .CLK(clk_bF_buf75), .D(_4917__3_), .Q(Ynonce_synth_3_) );
	DFFPOSX1 DFFPOSX1_382 ( .CLK(clk_bF_buf74), .D(_4917__4_), .Q(Ynonce_synth_4_) );
	DFFPOSX1 DFFPOSX1_383 ( .CLK(clk_bF_buf73), .D(_4917__5_), .Q(Ynonce_synth_5_) );
	DFFPOSX1 DFFPOSX1_384 ( .CLK(clk_bF_buf72), .D(_4917__6_), .Q(Ynonce_synth_6_) );
	DFFPOSX1 DFFPOSX1_385 ( .CLK(clk_bF_buf71), .D(_4917__7_), .Q(Ynonce_synth_7_) );
	DFFPOSX1 DFFPOSX1_386 ( .CLK(clk_bF_buf70), .D(_4917__8_), .Q(Ynonce_synth_8_) );
	DFFPOSX1 DFFPOSX1_387 ( .CLK(clk_bF_buf69), .D(_4917__9_), .Q(Ynonce_synth_9_) );
	DFFPOSX1 DFFPOSX1_388 ( .CLK(clk_bF_buf68), .D(_4917__10_), .Q(Ynonce_synth_10_) );
	DFFPOSX1 DFFPOSX1_389 ( .CLK(clk_bF_buf67), .D(_4917__11_), .Q(Ynonce_synth_11_) );
	DFFPOSX1 DFFPOSX1_390 ( .CLK(clk_bF_buf66), .D(_4917__12_), .Q(Ynonce_synth_12_) );
	DFFPOSX1 DFFPOSX1_391 ( .CLK(clk_bF_buf65), .D(_4917__13_), .Q(Ynonce_synth_13_) );
	DFFPOSX1 DFFPOSX1_392 ( .CLK(clk_bF_buf64), .D(_4917__14_), .Q(Ynonce_synth_14_) );
	DFFPOSX1 DFFPOSX1_393 ( .CLK(clk_bF_buf63), .D(_4917__15_), .Q(Ynonce_synth_15_) );
	DFFPOSX1 DFFPOSX1_394 ( .CLK(clk_bF_buf62), .D(_4917__16_), .Q(Ynonce_synth_16_) );
	DFFPOSX1 DFFPOSX1_395 ( .CLK(clk_bF_buf61), .D(_4917__17_), .Q(Ynonce_synth_17_) );
	DFFPOSX1 DFFPOSX1_396 ( .CLK(clk_bF_buf60), .D(_4917__18_), .Q(Ynonce_synth_18_) );
	DFFPOSX1 DFFPOSX1_397 ( .CLK(clk_bF_buf59), .D(_4917__19_), .Q(Ynonce_synth_19_) );
	DFFPOSX1 DFFPOSX1_398 ( .CLK(clk_bF_buf58), .D(_4917__20_), .Q(Ynonce_synth_20_) );
	DFFPOSX1 DFFPOSX1_399 ( .CLK(clk_bF_buf57), .D(_4917__21_), .Q(Ynonce_synth_21_) );
	DFFPOSX1 DFFPOSX1_400 ( .CLK(clk_bF_buf56), .D(_4917__22_), .Q(Ynonce_synth_22_) );
	DFFPOSX1 DFFPOSX1_401 ( .CLK(clk_bF_buf55), .D(_4917__23_), .Q(Ynonce_synth_23_) );
	DFFPOSX1 DFFPOSX1_402 ( .CLK(clk_bF_buf54), .D(_4917__24_), .Q(Ynonce_synth_24_) );
	DFFPOSX1 DFFPOSX1_403 ( .CLK(clk_bF_buf53), .D(_4917__25_), .Q(Ynonce_synth_25_) );
	DFFPOSX1 DFFPOSX1_404 ( .CLK(clk_bF_buf52), .D(_4917__26_), .Q(Ynonce_synth_26_) );
	DFFPOSX1 DFFPOSX1_405 ( .CLK(clk_bF_buf51), .D(_4917__27_), .Q(Ynonce_synth_27_) );
	DFFPOSX1 DFFPOSX1_406 ( .CLK(clk_bF_buf50), .D(_4917__28_), .Q(Ynonce_synth_28_) );
	DFFPOSX1 DFFPOSX1_407 ( .CLK(clk_bF_buf49), .D(_4917__29_), .Q(Ynonce_synth_29_) );
	DFFPOSX1 DFFPOSX1_408 ( .CLK(clk_bF_buf48), .D(_4917__30_), .Q(Ynonce_synth_30_) );
	DFFPOSX1 DFFPOSX1_409 ( .CLK(clk_bF_buf47), .D(_4917__31_), .Q(Ynonce_synth_31_) );
	DFFPOSX1 DFFPOSX1_410 ( .CLK(clk_bF_buf46), .D(_4918_), .Q(mux1_sel) );
	INVX8 INVX8_3 ( .A(reset_L_bF_buf0), .Y(_4997_) );
	INVX1 INVX1_283 ( .A(num_entradas[1]), .Y(_4998_) );
	INVX1 INVX1_284 ( .A(num_entradas[0]), .Y(_4999_) );
	OAI22X1 OAI22X1_208 ( .A(_4998_), .B(RAM_rd_ptr_1_), .C(_4999_), .D(RAM_rd_ptr_0_), .Y(_5000_) );
	INVX1 INVX1_285 ( .A(comparador_valid_bF_buf5), .Y(_5001_) );
	AOI21X1 AOI21X1_187 ( .A(RAM_rd_ptr_1_), .B(_4998_), .C(_5001_), .Y(_5002_) );
	AOI21X1 AOI21X1_188 ( .A(RAM_rd_ptr_0_), .B(_4999_), .C(_1__bF_buf5), .Y(_5003_) );
	OAI21X1 OAI21X1_391 ( .A(_5000_), .B(_5003_), .C(_5002_), .Y(_5004_) );
	NAND2X1 NAND2X1_192 ( .A(_3__0_), .B(_5004__bF_buf6), .Y(_5005_) );
	INVX1 INVX1_286 ( .A(RAM_rd_ptr_1_), .Y(_5006_) );
	INVX1 INVX1_287 ( .A(RAM_rd_ptr_0_), .Y(_5007_) );
	AOI22X1 AOI22X1_3 ( .A(_5006_), .B(num_entradas[1]), .C(num_entradas[0]), .D(_5007_), .Y(_5008_) );
	OAI21X1 OAI21X1_392 ( .A(_5006_), .B(num_entradas[1]), .C(comparador_valid_bF_buf4), .Y(_5009_) );
	INVX1 INVX1_288 ( .A(_1__bF_buf4), .Y(_5010_) );
	OAI21X1 OAI21X1_393 ( .A(_5007_), .B(num_entradas[0]), .C(_5010_), .Y(_5011_) );
	AOI21X1 AOI21X1_189 ( .A(_5011_), .B(_5008_), .C(_5009_), .Y(_5012_) );
	NAND2X1 NAND2X1_193 ( .A(comparador_nonce_synth_valido_0_), .B(_5012__bF_buf6), .Y(_5013_) );
	AOI21X1 AOI21X1_190 ( .A(_5005_), .B(_5013_), .C(_4997__bF_buf6), .Y(_4995__0_) );
	NAND2X1 NAND2X1_194 ( .A(_3__1_), .B(_5004__bF_buf5), .Y(_5014_) );
	NAND2X1 NAND2X1_195 ( .A(comparador_nonce_synth_valido_1_), .B(_5012__bF_buf5), .Y(_5015_) );
	AOI21X1 AOI21X1_191 ( .A(_5014_), .B(_5015_), .C(_4997__bF_buf5), .Y(_4995__1_) );
	NAND2X1 NAND2X1_196 ( .A(_3__2_), .B(_5004__bF_buf4), .Y(_5016_) );
	NAND2X1 NAND2X1_197 ( .A(comparador_nonce_synth_valido_2_), .B(_5012__bF_buf4), .Y(_5017_) );
	AOI21X1 AOI21X1_192 ( .A(_5016_), .B(_5017_), .C(_4997__bF_buf4), .Y(_4995__2_) );
	NAND2X1 NAND2X1_198 ( .A(_3__3_), .B(_5004__bF_buf3), .Y(_5018_) );
	NAND2X1 NAND2X1_199 ( .A(comparador_nonce_synth_valido_3_), .B(_5012__bF_buf3), .Y(_5019_) );
	AOI21X1 AOI21X1_193 ( .A(_5018_), .B(_5019_), .C(_4997__bF_buf3), .Y(_4995__3_) );
	NAND2X1 NAND2X1_200 ( .A(_3__4_), .B(_5004__bF_buf2), .Y(_5020_) );
	NAND2X1 NAND2X1_201 ( .A(comparador_nonce_synth_valido_4_), .B(_5012__bF_buf2), .Y(_5021_) );
	AOI21X1 AOI21X1_194 ( .A(_5020_), .B(_5021_), .C(_4997__bF_buf2), .Y(_4995__4_) );
	NAND2X1 NAND2X1_202 ( .A(_3__5_), .B(_5004__bF_buf1), .Y(_5022_) );
	NAND2X1 NAND2X1_203 ( .A(comparador_nonce_synth_valido_5_), .B(_5012__bF_buf1), .Y(_5023_) );
	AOI21X1 AOI21X1_195 ( .A(_5022_), .B(_5023_), .C(_4997__bF_buf1), .Y(_4995__5_) );
	NAND2X1 NAND2X1_204 ( .A(_3__6_), .B(_5004__bF_buf0), .Y(_5024_) );
	NAND2X1 NAND2X1_205 ( .A(comparador_nonce_synth_valido_6_), .B(_5012__bF_buf0), .Y(_5025_) );
	AOI21X1 AOI21X1_196 ( .A(_5024_), .B(_5025_), .C(_4997__bF_buf0), .Y(_4995__6_) );
	NAND2X1 NAND2X1_206 ( .A(_3__7_), .B(_5004__bF_buf6), .Y(_5026_) );
	NAND2X1 NAND2X1_207 ( .A(comparador_nonce_synth_valido_7_), .B(_5012__bF_buf6), .Y(_5027_) );
	AOI21X1 AOI21X1_197 ( .A(_5026_), .B(_5027_), .C(_4997__bF_buf6), .Y(_4995__7_) );
	NAND2X1 NAND2X1_208 ( .A(_3__8_), .B(_5004__bF_buf5), .Y(_5028_) );
	NAND2X1 NAND2X1_209 ( .A(comparador_nonce_synth_valido_8_), .B(_5012__bF_buf5), .Y(_5029_) );
	AOI21X1 AOI21X1_198 ( .A(_5028_), .B(_5029_), .C(_4997__bF_buf5), .Y(_4995__8_) );
	NAND2X1 NAND2X1_210 ( .A(_3__9_), .B(_5004__bF_buf4), .Y(_5030_) );
	NAND2X1 NAND2X1_211 ( .A(comparador_nonce_synth_valido_9_), .B(_5012__bF_buf4), .Y(_5031_) );
	AOI21X1 AOI21X1_199 ( .A(_5030_), .B(_5031_), .C(_4997__bF_buf4), .Y(_4995__9_) );
	NAND2X1 NAND2X1_212 ( .A(_3__10_), .B(_5004__bF_buf3), .Y(_5032_) );
	NAND2X1 NAND2X1_213 ( .A(comparador_nonce_synth_valido_10_), .B(_5012__bF_buf3), .Y(_5033_) );
	AOI21X1 AOI21X1_200 ( .A(_5032_), .B(_5033_), .C(_4997__bF_buf3), .Y(_4995__10_) );
	NAND2X1 NAND2X1_214 ( .A(_3__11_), .B(_5004__bF_buf2), .Y(_5034_) );
	NAND2X1 NAND2X1_215 ( .A(comparador_nonce_synth_valido_11_), .B(_5012__bF_buf2), .Y(_5035_) );
	AOI21X1 AOI21X1_201 ( .A(_5034_), .B(_5035_), .C(_4997__bF_buf2), .Y(_4995__11_) );
	NAND2X1 NAND2X1_216 ( .A(_3__12_), .B(_5004__bF_buf1), .Y(_5036_) );
	NAND2X1 NAND2X1_217 ( .A(comparador_nonce_synth_valido_12_), .B(_5012__bF_buf1), .Y(_5037_) );
	AOI21X1 AOI21X1_202 ( .A(_5036_), .B(_5037_), .C(_4997__bF_buf1), .Y(_4995__12_) );
	NAND2X1 NAND2X1_218 ( .A(_3__13_), .B(_5004__bF_buf0), .Y(_5038_) );
	NAND2X1 NAND2X1_219 ( .A(comparador_nonce_synth_valido_13_), .B(_5012__bF_buf0), .Y(_5039_) );
	AOI21X1 AOI21X1_203 ( .A(_5038_), .B(_5039_), .C(_4997__bF_buf0), .Y(_4995__13_) );
	NAND2X1 NAND2X1_220 ( .A(_3__14_), .B(_5004__bF_buf6), .Y(_5040_) );
	NAND2X1 NAND2X1_221 ( .A(comparador_nonce_synth_valido_14_), .B(_5012__bF_buf6), .Y(_5041_) );
	AOI21X1 AOI21X1_204 ( .A(_5040_), .B(_5041_), .C(_4997__bF_buf6), .Y(_4995__14_) );
	NAND2X1 NAND2X1_222 ( .A(_3__15_), .B(_5004__bF_buf5), .Y(_5042_) );
	NAND2X1 NAND2X1_223 ( .A(comparador_nonce_synth_valido_15_), .B(_5012__bF_buf5), .Y(_5043_) );
	AOI21X1 AOI21X1_205 ( .A(_5042_), .B(_5043_), .C(_4997__bF_buf5), .Y(_4995__15_) );
	NAND2X1 NAND2X1_224 ( .A(_3__16_), .B(_5004__bF_buf4), .Y(_5044_) );
	NAND2X1 NAND2X1_225 ( .A(comparador_nonce_synth_valido_16_), .B(_5012__bF_buf4), .Y(_5045_) );
	AOI21X1 AOI21X1_206 ( .A(_5044_), .B(_5045_), .C(_4997__bF_buf4), .Y(_4995__16_) );
	NAND2X1 NAND2X1_226 ( .A(_3__17_), .B(_5004__bF_buf3), .Y(_5046_) );
	NAND2X1 NAND2X1_227 ( .A(comparador_nonce_synth_valido_17_), .B(_5012__bF_buf3), .Y(_5047_) );
	AOI21X1 AOI21X1_207 ( .A(_5046_), .B(_5047_), .C(_4997__bF_buf3), .Y(_4995__17_) );
	NAND2X1 NAND2X1_228 ( .A(_3__18_), .B(_5004__bF_buf2), .Y(_5048_) );
	NAND2X1 NAND2X1_229 ( .A(comparador_nonce_synth_valido_18_), .B(_5012__bF_buf2), .Y(_5049_) );
	AOI21X1 AOI21X1_208 ( .A(_5048_), .B(_5049_), .C(_4997__bF_buf2), .Y(_4995__18_) );
	NAND2X1 NAND2X1_230 ( .A(_3__19_), .B(_5004__bF_buf1), .Y(_5050_) );
	NAND2X1 NAND2X1_231 ( .A(comparador_nonce_synth_valido_19_), .B(_5012__bF_buf1), .Y(_5051_) );
	AOI21X1 AOI21X1_209 ( .A(_5050_), .B(_5051_), .C(_4997__bF_buf1), .Y(_4995__19_) );
	NAND2X1 NAND2X1_232 ( .A(_3__20_), .B(_5004__bF_buf0), .Y(_5052_) );
	NAND2X1 NAND2X1_233 ( .A(comparador_nonce_synth_valido_20_), .B(_5012__bF_buf0), .Y(_5053_) );
	AOI21X1 AOI21X1_210 ( .A(_5052_), .B(_5053_), .C(_4997__bF_buf0), .Y(_4995__20_) );
	NAND2X1 NAND2X1_234 ( .A(_3__21_), .B(_5004__bF_buf6), .Y(_5054_) );
	NAND2X1 NAND2X1_235 ( .A(comparador_nonce_synth_valido_21_), .B(_5012__bF_buf6), .Y(_5055_) );
	AOI21X1 AOI21X1_211 ( .A(_5054_), .B(_5055_), .C(_4997__bF_buf6), .Y(_4995__21_) );
	NAND2X1 NAND2X1_236 ( .A(_3__22_), .B(_5004__bF_buf5), .Y(_5056_) );
	NAND2X1 NAND2X1_237 ( .A(comparador_nonce_synth_valido_22_), .B(_5012__bF_buf5), .Y(_5057_) );
	AOI21X1 AOI21X1_212 ( .A(_5056_), .B(_5057_), .C(_4997__bF_buf5), .Y(_4995__22_) );
	NAND2X1 NAND2X1_238 ( .A(_3__23_), .B(_5004__bF_buf4), .Y(_5058_) );
	NAND2X1 NAND2X1_239 ( .A(comparador_nonce_synth_valido_23_), .B(_5012__bF_buf4), .Y(_5059_) );
	AOI21X1 AOI21X1_213 ( .A(_5058_), .B(_5059_), .C(_4997__bF_buf4), .Y(_4995__23_) );
	NAND2X1 NAND2X1_240 ( .A(_3__24_), .B(_5004__bF_buf3), .Y(_5060_) );
	NAND2X1 NAND2X1_241 ( .A(comparador_nonce_synth_valido_24_), .B(_5012__bF_buf3), .Y(_5061_) );
	AOI21X1 AOI21X1_214 ( .A(_5060_), .B(_5061_), .C(_4997__bF_buf3), .Y(_4995__24_) );
	NAND2X1 NAND2X1_242 ( .A(_3__25_), .B(_5004__bF_buf2), .Y(_5062_) );
	NAND2X1 NAND2X1_243 ( .A(comparador_nonce_synth_valido_25_), .B(_5012__bF_buf2), .Y(_5063_) );
	AOI21X1 AOI21X1_215 ( .A(_5062_), .B(_5063_), .C(_4997__bF_buf2), .Y(_4995__25_) );
	NAND2X1 NAND2X1_244 ( .A(_3__26_), .B(_5004__bF_buf1), .Y(_5064_) );
	NAND2X1 NAND2X1_245 ( .A(comparador_nonce_synth_valido_26_), .B(_5012__bF_buf1), .Y(_5065_) );
	AOI21X1 AOI21X1_216 ( .A(_5064_), .B(_5065_), .C(_4997__bF_buf1), .Y(_4995__26_) );
	NAND2X1 NAND2X1_246 ( .A(_3__27_), .B(_5004__bF_buf0), .Y(_5066_) );
	NAND2X1 NAND2X1_247 ( .A(comparador_nonce_synth_valido_27_), .B(_5012__bF_buf0), .Y(_5067_) );
	AOI21X1 AOI21X1_217 ( .A(_5066_), .B(_5067_), .C(_4997__bF_buf0), .Y(_4995__27_) );
	NAND2X1 NAND2X1_248 ( .A(_3__28_), .B(_5004__bF_buf6), .Y(_5068_) );
	NAND2X1 NAND2X1_249 ( .A(comparador_nonce_synth_valido_28_), .B(_5012__bF_buf6), .Y(_5069_) );
	AOI21X1 AOI21X1_218 ( .A(_5068_), .B(_5069_), .C(_4997__bF_buf6), .Y(_4995__28_) );
	NAND2X1 NAND2X1_250 ( .A(_3__29_), .B(_5004__bF_buf5), .Y(_5070_) );
	NAND2X1 NAND2X1_251 ( .A(comparador_nonce_synth_valido_29_), .B(_5012__bF_buf5), .Y(_5071_) );
	AOI21X1 AOI21X1_219 ( .A(_5070_), .B(_5071_), .C(_4997__bF_buf5), .Y(_4995__29_) );
	NAND2X1 NAND2X1_252 ( .A(_3__30_), .B(_5004__bF_buf4), .Y(_5072_) );
	NAND2X1 NAND2X1_253 ( .A(comparador_nonce_synth_valido_30_), .B(_5012__bF_buf4), .Y(_5073_) );
	AOI21X1 AOI21X1_220 ( .A(_5072_), .B(_5073_), .C(_4997__bF_buf4), .Y(_4995__30_) );
	NAND2X1 NAND2X1_254 ( .A(_3__31_), .B(_5004__bF_buf3), .Y(_5074_) );
	NAND2X1 NAND2X1_255 ( .A(comparador_nonce_synth_valido_31_), .B(_5012__bF_buf3), .Y(_5075_) );
	AOI21X1 AOI21X1_221 ( .A(_5074_), .B(_5075_), .C(_4997__bF_buf3), .Y(_4995__31_) );
	NAND2X1 NAND2X1_256 ( .A(_0__0_), .B(_5004__bF_buf2), .Y(_5076_) );
	NAND2X1 NAND2X1_257 ( .A(bounty_synth_0_), .B(_5012__bF_buf2), .Y(_5077_) );
	AOI21X1 AOI21X1_222 ( .A(_5076_), .B(_5077_), .C(_4997__bF_buf2), .Y(_4993__0_) );
	NAND2X1 NAND2X1_258 ( .A(_0__1_), .B(_5004__bF_buf1), .Y(_5078_) );
	NAND2X1 NAND2X1_259 ( .A(bounty_synth_1_), .B(_5012__bF_buf1), .Y(_5079_) );
	AOI21X1 AOI21X1_223 ( .A(_5078_), .B(_5079_), .C(_4997__bF_buf1), .Y(_4993__1_) );
	NAND2X1 NAND2X1_260 ( .A(_0__2_), .B(_5004__bF_buf0), .Y(_5080_) );
	NAND2X1 NAND2X1_261 ( .A(bounty_synth_2_), .B(_5012__bF_buf0), .Y(_5081_) );
	AOI21X1 AOI21X1_224 ( .A(_5080_), .B(_5081_), .C(_4997__bF_buf0), .Y(_4993__2_) );
	NAND2X1 NAND2X1_262 ( .A(_0__3_), .B(_5004__bF_buf6), .Y(_5082_) );
	NAND2X1 NAND2X1_263 ( .A(bounty_synth_3_), .B(_5012__bF_buf6), .Y(_5083_) );
	AOI21X1 AOI21X1_225 ( .A(_5082_), .B(_5083_), .C(_4997__bF_buf6), .Y(_4993__3_) );
	NAND2X1 NAND2X1_264 ( .A(_0__4_), .B(_5004__bF_buf5), .Y(_5084_) );
	NAND2X1 NAND2X1_265 ( .A(bounty_synth_4_), .B(_5012__bF_buf5), .Y(_5085_) );
	AOI21X1 AOI21X1_226 ( .A(_5084_), .B(_5085_), .C(_4997__bF_buf5), .Y(_4993__4_) );
	NAND2X1 NAND2X1_266 ( .A(_0__5_), .B(_5004__bF_buf4), .Y(_5086_) );
	NAND2X1 NAND2X1_267 ( .A(bounty_synth_5_), .B(_5012__bF_buf4), .Y(_5087_) );
	AOI21X1 AOI21X1_227 ( .A(_5086_), .B(_5087_), .C(_4997__bF_buf4), .Y(_4993__5_) );
	NAND2X1 NAND2X1_268 ( .A(_0__6_), .B(_5004__bF_buf3), .Y(_5088_) );
	NAND2X1 NAND2X1_269 ( .A(bounty_synth_6_), .B(_5012__bF_buf3), .Y(_5089_) );
	AOI21X1 AOI21X1_228 ( .A(_5088_), .B(_5089_), .C(_4997__bF_buf3), .Y(_4993__6_) );
	NAND2X1 NAND2X1_270 ( .A(_0__7_), .B(_5004__bF_buf2), .Y(_5090_) );
	NAND2X1 NAND2X1_271 ( .A(bounty_synth_7_), .B(_5012__bF_buf2), .Y(_5091_) );
	AOI21X1 AOI21X1_229 ( .A(_5090_), .B(_5091_), .C(_4997__bF_buf2), .Y(_4993__7_) );
	NAND2X1 NAND2X1_272 ( .A(_0__8_), .B(_5004__bF_buf1), .Y(_5092_) );
	NAND2X1 NAND2X1_273 ( .A(bounty_synth_8_), .B(_5012__bF_buf1), .Y(_5093_) );
	AOI21X1 AOI21X1_230 ( .A(_5092_), .B(_5093_), .C(_4997__bF_buf1), .Y(_4993__8_) );
	NAND2X1 NAND2X1_274 ( .A(_0__9_), .B(_5004__bF_buf0), .Y(_5094_) );
	NAND2X1 NAND2X1_275 ( .A(bounty_synth_9_), .B(_5012__bF_buf0), .Y(_5095_) );
	AOI21X1 AOI21X1_231 ( .A(_5094_), .B(_5095_), .C(_4997__bF_buf0), .Y(_4993__9_) );
	NAND2X1 NAND2X1_276 ( .A(_0__10_), .B(_5004__bF_buf6), .Y(_5096_) );
	NAND2X1 NAND2X1_277 ( .A(bounty_synth_10_), .B(_5012__bF_buf6), .Y(_5097_) );
	AOI21X1 AOI21X1_232 ( .A(_5096_), .B(_5097_), .C(_4997__bF_buf6), .Y(_4993__10_) );
	NAND2X1 NAND2X1_278 ( .A(_0__11_), .B(_5004__bF_buf5), .Y(_5098_) );
	NAND2X1 NAND2X1_279 ( .A(bounty_synth_11_), .B(_5012__bF_buf5), .Y(_5099_) );
	AOI21X1 AOI21X1_233 ( .A(_5098_), .B(_5099_), .C(_4997__bF_buf5), .Y(_4993__11_) );
	NAND2X1 NAND2X1_280 ( .A(_0__12_), .B(_5004__bF_buf4), .Y(_5100_) );
	NAND2X1 NAND2X1_281 ( .A(bounty_synth_12_), .B(_5012__bF_buf4), .Y(_5101_) );
	AOI21X1 AOI21X1_234 ( .A(_5100_), .B(_5101_), .C(_4997__bF_buf4), .Y(_4993__12_) );
	NAND2X1 NAND2X1_282 ( .A(_0__13_), .B(_5004__bF_buf3), .Y(_5102_) );
	NAND2X1 NAND2X1_283 ( .A(bounty_synth_13_), .B(_5012__bF_buf3), .Y(_5103_) );
	AOI21X1 AOI21X1_235 ( .A(_5102_), .B(_5103_), .C(_4997__bF_buf3), .Y(_4993__13_) );
	NAND2X1 NAND2X1_284 ( .A(_0__14_), .B(_5004__bF_buf2), .Y(_5104_) );
	NAND2X1 NAND2X1_285 ( .A(bounty_synth_14_), .B(_5012__bF_buf2), .Y(_5105_) );
	AOI21X1 AOI21X1_236 ( .A(_5104_), .B(_5105_), .C(_4997__bF_buf2), .Y(_4993__14_) );
	NAND2X1 NAND2X1_286 ( .A(_0__15_), .B(_5004__bF_buf1), .Y(_5106_) );
	NAND2X1 NAND2X1_287 ( .A(bounty_synth_15_), .B(_5012__bF_buf1), .Y(_5107_) );
	AOI21X1 AOI21X1_237 ( .A(_5106_), .B(_5107_), .C(_4997__bF_buf1), .Y(_4993__15_) );
	NAND2X1 NAND2X1_288 ( .A(_0__16_), .B(_5004__bF_buf0), .Y(_5108_) );
	NAND2X1 NAND2X1_289 ( .A(bounty_synth_16_), .B(_5012__bF_buf0), .Y(_5109_) );
	AOI21X1 AOI21X1_238 ( .A(_5108_), .B(_5109_), .C(_4997__bF_buf0), .Y(_4993__16_) );
	NAND2X1 NAND2X1_290 ( .A(_0__17_), .B(_5004__bF_buf6), .Y(_5110_) );
	NAND2X1 NAND2X1_291 ( .A(bounty_synth_17_), .B(_5012__bF_buf6), .Y(_5111_) );
	AOI21X1 AOI21X1_239 ( .A(_5110_), .B(_5111_), .C(_4997__bF_buf6), .Y(_4993__17_) );
	NAND2X1 NAND2X1_292 ( .A(_0__18_), .B(_5004__bF_buf5), .Y(_5112_) );
	NAND2X1 NAND2X1_293 ( .A(bounty_synth_18_), .B(_5012__bF_buf5), .Y(_5113_) );
	AOI21X1 AOI21X1_240 ( .A(_5112_), .B(_5113_), .C(_4997__bF_buf5), .Y(_4993__18_) );
	NAND2X1 NAND2X1_294 ( .A(_0__19_), .B(_5004__bF_buf4), .Y(_5114_) );
	NAND2X1 NAND2X1_295 ( .A(bounty_synth_19_), .B(_5012__bF_buf4), .Y(_5115_) );
	AOI21X1 AOI21X1_241 ( .A(_5114_), .B(_5115_), .C(_4997__bF_buf4), .Y(_4993__19_) );
	NAND2X1 NAND2X1_296 ( .A(_0__20_), .B(_5004__bF_buf3), .Y(_5116_) );
	NAND2X1 NAND2X1_297 ( .A(bounty_synth_20_), .B(_5012__bF_buf3), .Y(_5117_) );
	AOI21X1 AOI21X1_242 ( .A(_5116_), .B(_5117_), .C(_4997__bF_buf3), .Y(_4993__20_) );
	NAND2X1 NAND2X1_298 ( .A(_0__21_), .B(_5004__bF_buf2), .Y(_5118_) );
	NAND2X1 NAND2X1_299 ( .A(bounty_synth_21_), .B(_5012__bF_buf2), .Y(_5119_) );
	AOI21X1 AOI21X1_243 ( .A(_5118_), .B(_5119_), .C(_4997__bF_buf2), .Y(_4993__21_) );
	NAND2X1 NAND2X1_300 ( .A(_0__22_), .B(_5004__bF_buf1), .Y(_5120_) );
	NAND2X1 NAND2X1_301 ( .A(bounty_synth_22_), .B(_5012__bF_buf1), .Y(_5121_) );
	AOI21X1 AOI21X1_244 ( .A(_5120_), .B(_5121_), .C(_4997__bF_buf1), .Y(_4993__22_) );
	NAND2X1 NAND2X1_302 ( .A(_0__23_), .B(_5004__bF_buf0), .Y(_5122_) );
	NAND2X1 NAND2X1_303 ( .A(bounty_synth_23_), .B(_5012__bF_buf0), .Y(_5123_) );
	AOI21X1 AOI21X1_245 ( .A(_5122_), .B(_5123_), .C(_4997__bF_buf0), .Y(_4993__23_) );
	OAI21X1 OAI21X1_394 ( .A(_5008_), .B(_5009_), .C(RAM_rd_ptr_0_), .Y(_5124_) );
	NAND3X1 NAND3X1_58 ( .A(_5007_), .B(_5002_), .C(_5000_), .Y(_5125_) );
	AOI21X1 AOI21X1_246 ( .A(_5125_), .B(_5124_), .C(_4997__bF_buf6), .Y(_4996__0_) );
	NAND3X1 NAND3X1_59 ( .A(num_entradas[1]), .B(RAM_rd_ptr_0_), .C(comparador_valid_bF_buf3), .Y(_5126_) );
	AOI21X1 AOI21X1_247 ( .A(_5006_), .B(_5126_), .C(_4997__bF_buf5), .Y(_4996__1_) );
	NAND3X1 NAND3X1_60 ( .A(_5002_), .B(_5003_), .C(_5008_), .Y(_5127_) );
	OAI21X1 OAI21X1_395 ( .A(_5008_), .B(_5009_), .C(_1__bF_buf3), .Y(_5128_) );
	AOI21X1 AOI21X1_248 ( .A(_5127_), .B(_5128_), .C(_4997__bF_buf4), .Y(_4994_) );
	DFFPOSX1 DFFPOSX1_411 ( .CLK(clk_bF_buf45), .D(_4994_), .Q(_1_) );
	DFFPOSX1 DFFPOSX1_412 ( .CLK(clk_bF_buf44), .D(_4996__0_), .Q(RAM_rd_ptr_0_) );
	DFFPOSX1 DFFPOSX1_413 ( .CLK(clk_bF_buf43), .D(_4996__1_), .Q(RAM_rd_ptr_1_) );
	DFFPOSX1 DFFPOSX1_414 ( .CLK(clk_bF_buf42), .D(_4993__0_), .Q(_0__0_) );
	DFFPOSX1 DFFPOSX1_415 ( .CLK(clk_bF_buf41), .D(_4993__1_), .Q(_0__1_) );
	DFFPOSX1 DFFPOSX1_416 ( .CLK(clk_bF_buf40), .D(_4993__2_), .Q(_0__2_) );
	DFFPOSX1 DFFPOSX1_417 ( .CLK(clk_bF_buf39), .D(_4993__3_), .Q(_0__3_) );
	DFFPOSX1 DFFPOSX1_418 ( .CLK(clk_bF_buf38), .D(_4993__4_), .Q(_0__4_) );
	DFFPOSX1 DFFPOSX1_419 ( .CLK(clk_bF_buf37), .D(_4993__5_), .Q(_0__5_) );
	DFFPOSX1 DFFPOSX1_420 ( .CLK(clk_bF_buf36), .D(_4993__6_), .Q(_0__6_) );
	DFFPOSX1 DFFPOSX1_421 ( .CLK(clk_bF_buf35), .D(_4993__7_), .Q(_0__7_) );
	DFFPOSX1 DFFPOSX1_422 ( .CLK(clk_bF_buf34), .D(_4993__8_), .Q(_0__8_) );
	DFFPOSX1 DFFPOSX1_423 ( .CLK(clk_bF_buf33), .D(_4993__9_), .Q(_0__9_) );
	DFFPOSX1 DFFPOSX1_424 ( .CLK(clk_bF_buf32), .D(_4993__10_), .Q(_0__10_) );
	DFFPOSX1 DFFPOSX1_425 ( .CLK(clk_bF_buf31), .D(_4993__11_), .Q(_0__11_) );
	DFFPOSX1 DFFPOSX1_426 ( .CLK(clk_bF_buf30), .D(_4993__12_), .Q(_0__12_) );
	DFFPOSX1 DFFPOSX1_427 ( .CLK(clk_bF_buf29), .D(_4993__13_), .Q(_0__13_) );
	DFFPOSX1 DFFPOSX1_428 ( .CLK(clk_bF_buf28), .D(_4993__14_), .Q(_0__14_) );
	DFFPOSX1 DFFPOSX1_429 ( .CLK(clk_bF_buf27), .D(_4993__15_), .Q(_0__15_) );
	DFFPOSX1 DFFPOSX1_430 ( .CLK(clk_bF_buf26), .D(_4993__16_), .Q(_0__16_) );
	DFFPOSX1 DFFPOSX1_431 ( .CLK(clk_bF_buf25), .D(_4993__17_), .Q(_0__17_) );
	DFFPOSX1 DFFPOSX1_432 ( .CLK(clk_bF_buf24), .D(_4993__18_), .Q(_0__18_) );
	DFFPOSX1 DFFPOSX1_433 ( .CLK(clk_bF_buf23), .D(_4993__19_), .Q(_0__19_) );
	DFFPOSX1 DFFPOSX1_434 ( .CLK(clk_bF_buf22), .D(_4993__20_), .Q(_0__20_) );
	DFFPOSX1 DFFPOSX1_435 ( .CLK(clk_bF_buf21), .D(_4993__21_), .Q(_0__21_) );
	DFFPOSX1 DFFPOSX1_436 ( .CLK(clk_bF_buf20), .D(_4993__22_), .Q(_0__22_) );
	DFFPOSX1 DFFPOSX1_437 ( .CLK(clk_bF_buf19), .D(_4993__23_), .Q(_0__23_) );
	DFFPOSX1 DFFPOSX1_438 ( .CLK(clk_bF_buf18), .D(_4995__0_), .Q(_3__0_) );
	DFFPOSX1 DFFPOSX1_439 ( .CLK(clk_bF_buf17), .D(_4995__1_), .Q(_3__1_) );
	DFFPOSX1 DFFPOSX1_440 ( .CLK(clk_bF_buf16), .D(_4995__2_), .Q(_3__2_) );
	DFFPOSX1 DFFPOSX1_441 ( .CLK(clk_bF_buf15), .D(_4995__3_), .Q(_3__3_) );
	DFFPOSX1 DFFPOSX1_442 ( .CLK(clk_bF_buf14), .D(_4995__4_), .Q(_3__4_) );
	DFFPOSX1 DFFPOSX1_443 ( .CLK(clk_bF_buf13), .D(_4995__5_), .Q(_3__5_) );
	DFFPOSX1 DFFPOSX1_444 ( .CLK(clk_bF_buf12), .D(_4995__6_), .Q(_3__6_) );
	DFFPOSX1 DFFPOSX1_445 ( .CLK(clk_bF_buf11), .D(_4995__7_), .Q(_3__7_) );
	DFFPOSX1 DFFPOSX1_446 ( .CLK(clk_bF_buf10), .D(_4995__8_), .Q(_3__8_) );
	DFFPOSX1 DFFPOSX1_447 ( .CLK(clk_bF_buf9), .D(_4995__9_), .Q(_3__9_) );
	DFFPOSX1 DFFPOSX1_448 ( .CLK(clk_bF_buf8), .D(_4995__10_), .Q(_3__10_) );
	DFFPOSX1 DFFPOSX1_449 ( .CLK(clk_bF_buf7), .D(_4995__11_), .Q(_3__11_) );
	DFFPOSX1 DFFPOSX1_450 ( .CLK(clk_bF_buf6), .D(_4995__12_), .Q(_3__12_) );
	DFFPOSX1 DFFPOSX1_451 ( .CLK(clk_bF_buf5), .D(_4995__13_), .Q(_3__13_) );
	DFFPOSX1 DFFPOSX1_452 ( .CLK(clk_bF_buf4), .D(_4995__14_), .Q(_3__14_) );
	DFFPOSX1 DFFPOSX1_453 ( .CLK(clk_bF_buf3), .D(_4995__15_), .Q(_3__15_) );
	DFFPOSX1 DFFPOSX1_454 ( .CLK(clk_bF_buf2), .D(_4995__16_), .Q(_3__16_) );
	DFFPOSX1 DFFPOSX1_455 ( .CLK(clk_bF_buf1), .D(_4995__17_), .Q(_3__17_) );
	DFFPOSX1 DFFPOSX1_456 ( .CLK(clk_bF_buf0), .D(_4995__18_), .Q(_3__18_) );
	DFFPOSX1 DFFPOSX1_457 ( .CLK(clk_bF_buf113), .D(_4995__19_), .Q(_3__19_) );
	DFFPOSX1 DFFPOSX1_458 ( .CLK(clk_bF_buf112), .D(_4995__20_), .Q(_3__20_) );
	DFFPOSX1 DFFPOSX1_459 ( .CLK(clk_bF_buf111), .D(_4995__21_), .Q(_3__21_) );
	DFFPOSX1 DFFPOSX1_460 ( .CLK(clk_bF_buf110), .D(_4995__22_), .Q(_3__22_) );
	DFFPOSX1 DFFPOSX1_461 ( .CLK(clk_bF_buf109), .D(_4995__23_), .Q(_3__23_) );
	DFFPOSX1 DFFPOSX1_462 ( .CLK(clk_bF_buf108), .D(_4995__24_), .Q(_3__24_) );
	DFFPOSX1 DFFPOSX1_463 ( .CLK(clk_bF_buf107), .D(_4995__25_), .Q(_3__25_) );
	DFFPOSX1 DFFPOSX1_464 ( .CLK(clk_bF_buf106), .D(_4995__26_), .Q(_3__26_) );
	DFFPOSX1 DFFPOSX1_465 ( .CLK(clk_bF_buf105), .D(_4995__27_), .Q(_3__27_) );
	DFFPOSX1 DFFPOSX1_466 ( .CLK(clk_bF_buf104), .D(_4995__28_), .Q(_3__28_) );
	DFFPOSX1 DFFPOSX1_467 ( .CLK(clk_bF_buf103), .D(_4995__29_), .Q(_3__29_) );
	DFFPOSX1 DFFPOSX1_468 ( .CLK(clk_bF_buf102), .D(_4995__30_), .Q(_3__30_) );
	DFFPOSX1 DFFPOSX1_469 ( .CLK(clk_bF_buf101), .D(_4995__31_), .Q(_3__31_) );
	BUFX2 BUFX2_279 ( .A(_0__0_), .Y(bounty_synth_out[0]) );
	BUFX2 BUFX2_280 ( .A(_0__1_), .Y(bounty_synth_out[1]) );
	BUFX2 BUFX2_281 ( .A(_0__2_), .Y(bounty_synth_out[2]) );
	BUFX2 BUFX2_282 ( .A(_0__3_), .Y(bounty_synth_out[3]) );
	BUFX2 BUFX2_283 ( .A(_0__4_), .Y(bounty_synth_out[4]) );
	BUFX2 BUFX2_284 ( .A(_0__5_), .Y(bounty_synth_out[5]) );
	BUFX2 BUFX2_285 ( .A(_0__6_), .Y(bounty_synth_out[6]) );
	BUFX2 BUFX2_286 ( .A(_0__7_), .Y(bounty_synth_out[7]) );
	BUFX2 BUFX2_287 ( .A(_0__8_), .Y(bounty_synth_out[8]) );
	BUFX2 BUFX2_288 ( .A(_0__9_), .Y(bounty_synth_out[9]) );
	BUFX2 BUFX2_289 ( .A(_0__10_), .Y(bounty_synth_out[10]) );
	BUFX2 BUFX2_290 ( .A(_0__11_), .Y(bounty_synth_out[11]) );
	BUFX2 BUFX2_291 ( .A(_0__12_), .Y(bounty_synth_out[12]) );
	BUFX2 BUFX2_292 ( .A(_0__13_), .Y(bounty_synth_out[13]) );
	BUFX2 BUFX2_293 ( .A(_0__14_), .Y(bounty_synth_out[14]) );
	BUFX2 BUFX2_294 ( .A(_0__15_), .Y(bounty_synth_out[15]) );
	BUFX2 BUFX2_295 ( .A(_0__16_), .Y(bounty_synth_out[16]) );
	BUFX2 BUFX2_296 ( .A(_0__17_), .Y(bounty_synth_out[17]) );
	BUFX2 BUFX2_297 ( .A(_0__18_), .Y(bounty_synth_out[18]) );
	BUFX2 BUFX2_298 ( .A(_0__19_), .Y(bounty_synth_out[19]) );
	BUFX2 BUFX2_299 ( .A(_0__20_), .Y(bounty_synth_out[20]) );
	BUFX2 BUFX2_300 ( .A(_0__21_), .Y(bounty_synth_out[21]) );
	BUFX2 BUFX2_301 ( .A(_0__22_), .Y(bounty_synth_out[22]) );
	BUFX2 BUFX2_302 ( .A(_0__23_), .Y(bounty_synth_out[23]) );
	BUFX2 BUFX2_303 ( .A(_1__bF_buf2), .Y(fin_synth) );
	BUFX2 BUFX2_304 ( .A(_2__0_), .Y(nonce_synth[0]) );
	BUFX2 BUFX2_305 ( .A(_2__1_), .Y(nonce_synth[1]) );
	BUFX2 BUFX2_306 ( .A(_2__2_), .Y(nonce_synth[2]) );
	BUFX2 BUFX2_307 ( .A(_2__3_), .Y(nonce_synth[3]) );
	BUFX2 BUFX2_308 ( .A(_2__4_), .Y(nonce_synth[4]) );
	BUFX2 BUFX2_309 ( .A(_2__5_), .Y(nonce_synth[5]) );
	BUFX2 BUFX2_310 ( .A(_2__6_), .Y(nonce_synth[6]) );
	BUFX2 BUFX2_311 ( .A(_2__7_), .Y(nonce_synth[7]) );
	BUFX2 BUFX2_312 ( .A(_2__8_), .Y(nonce_synth[8]) );
	BUFX2 BUFX2_313 ( .A(_2__9_), .Y(nonce_synth[9]) );
	BUFX2 BUFX2_314 ( .A(_2__10_), .Y(nonce_synth[10]) );
	BUFX2 BUFX2_315 ( .A(_2__11_), .Y(nonce_synth[11]) );
	BUFX2 BUFX2_316 ( .A(_2__12_), .Y(nonce_synth[12]) );
	BUFX2 BUFX2_317 ( .A(_2__13_), .Y(nonce_synth[13]) );
	BUFX2 BUFX2_318 ( .A(_2__14_), .Y(nonce_synth[14]) );
	BUFX2 BUFX2_319 ( .A(_2__15_), .Y(nonce_synth[15]) );
	BUFX2 BUFX2_320 ( .A(_2__16_), .Y(nonce_synth[16]) );
	BUFX2 BUFX2_321 ( .A(_2__17_), .Y(nonce_synth[17]) );
	BUFX2 BUFX2_322 ( .A(_2__18_), .Y(nonce_synth[18]) );
	BUFX2 BUFX2_323 ( .A(_2__19_), .Y(nonce_synth[19]) );
	BUFX2 BUFX2_324 ( .A(_2__20_), .Y(nonce_synth[20]) );
	BUFX2 BUFX2_325 ( .A(_2__21_), .Y(nonce_synth[21]) );
	BUFX2 BUFX2_326 ( .A(_2__22_), .Y(nonce_synth[22]) );
	BUFX2 BUFX2_327 ( .A(_2__23_), .Y(nonce_synth[23]) );
	BUFX2 BUFX2_328 ( .A(_2__24_), .Y(nonce_synth[24]) );
	BUFX2 BUFX2_329 ( .A(_2__25_), .Y(nonce_synth[25]) );
	BUFX2 BUFX2_330 ( .A(_2__26_), .Y(nonce_synth[26]) );
	BUFX2 BUFX2_331 ( .A(_2__27_), .Y(nonce_synth[27]) );
	BUFX2 BUFX2_332 ( .A(_2__28_), .Y(nonce_synth[28]) );
	BUFX2 BUFX2_333 ( .A(_2__29_), .Y(nonce_synth[29]) );
	BUFX2 BUFX2_334 ( .A(_2__30_), .Y(nonce_synth[30]) );
	BUFX2 BUFX2_335 ( .A(_2__31_), .Y(nonce_synth[31]) );
	BUFX2 BUFX2_336 ( .A(_3__0_), .Y(nonce_synth_valido_out[0]) );
	BUFX2 BUFX2_337 ( .A(_3__1_), .Y(nonce_synth_valido_out[1]) );
	BUFX2 BUFX2_338 ( .A(_3__2_), .Y(nonce_synth_valido_out[2]) );
	BUFX2 BUFX2_339 ( .A(_3__3_), .Y(nonce_synth_valido_out[3]) );
	BUFX2 BUFX2_340 ( .A(_3__4_), .Y(nonce_synth_valido_out[4]) );
	BUFX2 BUFX2_341 ( .A(_3__5_), .Y(nonce_synth_valido_out[5]) );
	BUFX2 BUFX2_342 ( .A(_3__6_), .Y(nonce_synth_valido_out[6]) );
	BUFX2 BUFX2_343 ( .A(_3__7_), .Y(nonce_synth_valido_out[7]) );
	BUFX2 BUFX2_344 ( .A(_3__8_), .Y(nonce_synth_valido_out[8]) );
	BUFX2 BUFX2_345 ( .A(_3__9_), .Y(nonce_synth_valido_out[9]) );
	BUFX2 BUFX2_346 ( .A(_3__10_), .Y(nonce_synth_valido_out[10]) );
	BUFX2 BUFX2_347 ( .A(_3__11_), .Y(nonce_synth_valido_out[11]) );
	BUFX2 BUFX2_348 ( .A(_3__12_), .Y(nonce_synth_valido_out[12]) );
	BUFX2 BUFX2_349 ( .A(_3__13_), .Y(nonce_synth_valido_out[13]) );
	BUFX2 BUFX2_350 ( .A(_3__14_), .Y(nonce_synth_valido_out[14]) );
	BUFX2 BUFX2_351 ( .A(_3__15_), .Y(nonce_synth_valido_out[15]) );
	BUFX2 BUFX2_352 ( .A(_3__16_), .Y(nonce_synth_valido_out[16]) );
	BUFX2 BUFX2_353 ( .A(_3__17_), .Y(nonce_synth_valido_out[17]) );
	BUFX2 BUFX2_354 ( .A(_3__18_), .Y(nonce_synth_valido_out[18]) );
	BUFX2 BUFX2_355 ( .A(_3__19_), .Y(nonce_synth_valido_out[19]) );
	BUFX2 BUFX2_356 ( .A(_3__20_), .Y(nonce_synth_valido_out[20]) );
	BUFX2 BUFX2_357 ( .A(_3__21_), .Y(nonce_synth_valido_out[21]) );
	BUFX2 BUFX2_358 ( .A(_3__22_), .Y(nonce_synth_valido_out[22]) );
	BUFX2 BUFX2_359 ( .A(_3__23_), .Y(nonce_synth_valido_out[23]) );
	BUFX2 BUFX2_360 ( .A(_3__24_), .Y(nonce_synth_valido_out[24]) );
	BUFX2 BUFX2_361 ( .A(_3__25_), .Y(nonce_synth_valido_out[25]) );
	BUFX2 BUFX2_362 ( .A(_3__26_), .Y(nonce_synth_valido_out[26]) );
	BUFX2 BUFX2_363 ( .A(_3__27_), .Y(nonce_synth_valido_out[27]) );
	BUFX2 BUFX2_364 ( .A(_3__28_), .Y(nonce_synth_valido_out[28]) );
	BUFX2 BUFX2_365 ( .A(_3__29_), .Y(nonce_synth_valido_out[29]) );
	BUFX2 BUFX2_366 ( .A(_3__30_), .Y(nonce_synth_valido_out[30]) );
	BUFX2 BUFX2_367 ( .A(_3__31_), .Y(nonce_synth_valido_out[31]) );
	NAND2X1 NAND2X1_304 ( .A(reset_L_bF_buf49), .B(RAM_rd_ptr_0_), .Y(_4__88_) );
	INVX1 INVX1_289 ( .A(_4__88_), .Y(_4__89_) );
	NAND2X1 NAND2X1_305 ( .A(reset_L_bF_buf48), .B(RAM_rd_ptr_1_), .Y(_4__92_) );
	INVX1 INVX1_290 ( .A(_4__92_), .Y(_4__77_) );
	OR2X2 OR2X2_16 ( .A(_4__88_), .B(RAM_rd_ptr_1_), .Y(_4__84_) );
	NOR2X1 NOR2X1_188 ( .A(RAM_rd_ptr_0_), .B(_4__92_), .Y(_4__94_) );
	NAND3X1 NAND3X1_61 ( .A(reset_L_bF_buf47), .B(RAM_rd_ptr_0_), .C(RAM_rd_ptr_1_), .Y(_4__93_) );
	OAI21X1 OAI21X1_396 ( .A(RAM_rd_ptr_0_), .B(RAM_rd_ptr_1_), .C(reset_L_bF_buf46), .Y(_4__82_) );
	INVX1 INVX1_291 ( .A(_4__82_), .Y(_4__95_) );
	NAND2X1 NAND2X1_306 ( .A(RAM_rd_ptr_0_), .B(RAM_rd_ptr_1_), .Y(_5_) );
	OR2X2 OR2X2_17 ( .A(RAM_rd_ptr_0_), .B(RAM_rd_ptr_1_), .Y(_6_) );
	NAND3X1 NAND3X1_62 ( .A(reset_L_bF_buf45), .B(_5_), .C(_6_), .Y(_4__86_) );
	AOI21X1 AOI21X1_249 ( .A(RAM_rd_ptr_0_), .B(RAM_rd_ptr_1_), .C(_4__82_), .Y(_4__46_) );
	INVX1 INVX1_292 ( .A(_4__93_), .Y(_4__71_) );
	NOR2X1 NOR2X1_189 ( .A(RAM_rd_ptr_1_), .B(_4__88_), .Y(_4__58_) );
	OR2X2 OR2X2_18 ( .A(_4__92_), .B(RAM_rd_ptr_0_), .Y(_4__85_) );
	DFFPOSX1 DFFPOSX1_470 ( .CLK(clk_bF_buf100), .D(_4__46_), .Q(RAM_entrada_46_) );
	DFFPOSX1 DFFPOSX1_471 ( .CLK(clk_bF_buf99), .D(_4__58_), .Q(RAM_entrada_58_) );
	DFFPOSX1 DFFPOSX1_472 ( .CLK(clk_bF_buf98), .D(_4__95_), .Q(RAM_entrada_95_) );
	DFFPOSX1 DFFPOSX1_473 ( .CLK(clk_bF_buf97), .D(_4__71_), .Q(RAM_entrada_71_) );
	DFFPOSX1 DFFPOSX1_474 ( .CLK(clk_bF_buf96), .D(_4__77_), .Q(RAM_entrada_77_) );
	DFFPOSX1 DFFPOSX1_475 ( .CLK(clk_bF_buf95), .D(_4__82_), .Q(RAM_entrada_82_) );
	DFFPOSX1 DFFPOSX1_476 ( .CLK(clk_bF_buf94), .D(_4__84_), .Q(RAM_entrada_84_) );
	DFFPOSX1 DFFPOSX1_477 ( .CLK(clk_bF_buf93), .D(_4__85_), .Q(RAM_entrada_85_) );
	DFFPOSX1 DFFPOSX1_478 ( .CLK(clk_bF_buf92), .D(_4__86_), .Q(RAM_entrada_86_) );
	DFFPOSX1 DFFPOSX1_479 ( .CLK(clk_bF_buf91), .D(_4__88_), .Q(RAM_entrada_88_) );
	DFFPOSX1 DFFPOSX1_480 ( .CLK(clk_bF_buf90), .D(_4__89_), .Q(RAM_entrada_89_) );
	DFFPOSX1 DFFPOSX1_481 ( .CLK(clk_bF_buf89), .D(_4__92_), .Q(RAM_entrada_92_) );
	DFFPOSX1 DFFPOSX1_482 ( .CLK(clk_bF_buf88), .D(_4__93_), .Q(RAM_entrada_93_) );
	DFFPOSX1 DFFPOSX1_483 ( .CLK(clk_bF_buf87), .D(_4__94_), .Q(RAM_entrada_94_) );
	INVX8 INVX8_4 ( .A(reset_L_bF_buf44), .Y(_10_) );
	INVX1 INVX1_293 ( .A(Y_17_), .Y(_11_) );
	NOR2X1 NOR2X1_190 ( .A(target[1]), .B(_11_), .Y(_12_) );
	INVX1 INVX1_294 ( .A(Y_16_), .Y(_13_) );
	NAND2X1 NAND2X1_307 ( .A(target[0]), .B(_13_), .Y(_14_) );
	NAND2X1 NAND2X1_308 ( .A(target[1]), .B(_11_), .Y(_15_) );
	AOI21X1 AOI21X1_250 ( .A(_14_), .B(_15_), .C(_12_), .Y(_16_) );
	AND2X2 AND2X2_32 ( .A(target[3]), .B(Y_19_), .Y(_17_) );
	NOR2X1 NOR2X1_191 ( .A(target[3]), .B(Y_19_), .Y(_18_) );
	NAND2X1 NAND2X1_309 ( .A(target[2]), .B(Y_18_), .Y(_19_) );
	INVX1 INVX1_295 ( .A(_19_), .Y(_20_) );
	NOR2X1 NOR2X1_192 ( .A(target[2]), .B(Y_18_), .Y(_21_) );
	OAI22X1 OAI22X1_209 ( .A(_17_), .B(_18_), .C(_20_), .D(_21_), .Y(_22_) );
	INVX1 INVX1_296 ( .A(Y_19_), .Y(_23_) );
	NOR2X1 NOR2X1_193 ( .A(target[3]), .B(_23_), .Y(_24_) );
	NAND2X1 NAND2X1_310 ( .A(target[3]), .B(_23_), .Y(_25_) );
	INVX1 INVX1_297 ( .A(Y_18_), .Y(_26_) );
	NOR2X1 NOR2X1_194 ( .A(target[2]), .B(_26_), .Y(_27_) );
	AOI21X1 AOI21X1_251 ( .A(_25_), .B(_27_), .C(_24_), .Y(_28_) );
	OAI21X1 OAI21X1_397 ( .A(_22_), .B(_16_), .C(_28_), .Y(_29_) );
	NAND2X1 NAND2X1_311 ( .A(target[7]), .B(Y_23_), .Y(_30_) );
	INVX1 INVX1_298 ( .A(_30_), .Y(_31_) );
	NOR2X1 NOR2X1_195 ( .A(target[7]), .B(Y_23_), .Y(_32_) );
	NAND2X1 NAND2X1_312 ( .A(target[6]), .B(Y_22_), .Y(_33_) );
	INVX1 INVX1_299 ( .A(_33_), .Y(_34_) );
	NOR2X1 NOR2X1_196 ( .A(target[6]), .B(Y_22_), .Y(_35_) );
	OAI22X1 OAI22X1_210 ( .A(_31_), .B(_32_), .C(_34_), .D(_35_), .Y(_36_) );
	INVX1 INVX1_300 ( .A(target[5]), .Y(_37_) );
	INVX1 INVX1_301 ( .A(target[4]), .Y(_38_) );
	AOI22X1 AOI22X1_4 ( .A(_37_), .B(Y_21_), .C(_38_), .D(Y_20_), .Y(_39_) );
	INVX1 INVX1_302 ( .A(Y_21_), .Y(_40_) );
	INVX1 INVX1_303 ( .A(Y_20_), .Y(_41_) );
	AOI22X1 AOI22X1_5 ( .A(_40_), .B(target[5]), .C(target[4]), .D(_41_), .Y(_42_) );
	NAND2X1 NAND2X1_313 ( .A(_39_), .B(_42_), .Y(_43_) );
	NOR2X1 NOR2X1_197 ( .A(_36_), .B(_43_), .Y(_44_) );
	INVX1 INVX1_304 ( .A(target[7]), .Y(_45_) );
	INVX1 INVX1_305 ( .A(Y_23_), .Y(_46_) );
	INVX1 INVX1_306 ( .A(Y_22_), .Y(_47_) );
	OAI22X1 OAI22X1_211 ( .A(_46_), .B(target[7]), .C(target[6]), .D(_47_), .Y(_48_) );
	OAI21X1 OAI21X1_398 ( .A(_45_), .B(Y_23_), .C(_48_), .Y(_49_) );
	OAI22X1 OAI22X1_212 ( .A(_40_), .B(target[5]), .C(target[4]), .D(_41_), .Y(_50_) );
	OAI21X1 OAI21X1_399 ( .A(_37_), .B(Y_21_), .C(_50_), .Y(_51_) );
	OAI21X1 OAI21X1_400 ( .A(_51_), .B(_36_), .C(_49_), .Y(_52_) );
	AOI21X1 AOI21X1_252 ( .A(_44_), .B(_29_), .C(_52_), .Y(_53_) );
	INVX1 INVX1_307 ( .A(Y_9_), .Y(_54_) );
	NOR2X1 NOR2X1_198 ( .A(target[1]), .B(_54_), .Y(_55_) );
	INVX1 INVX1_308 ( .A(Y_8_), .Y(_56_) );
	NAND2X1 NAND2X1_314 ( .A(target[0]), .B(_56_), .Y(_57_) );
	NAND2X1 NAND2X1_315 ( .A(target[1]), .B(_54_), .Y(_58_) );
	AOI21X1 AOI21X1_253 ( .A(_57_), .B(_58_), .C(_55_), .Y(_59_) );
	NAND2X1 NAND2X1_316 ( .A(target[3]), .B(Y_11_), .Y(_60_) );
	INVX1 INVX1_309 ( .A(_60_), .Y(_61_) );
	NOR2X1 NOR2X1_199 ( .A(target[3]), .B(Y_11_), .Y(_62_) );
	NAND2X1 NAND2X1_317 ( .A(target[2]), .B(Y_10_), .Y(_63_) );
	INVX1 INVX1_310 ( .A(_63_), .Y(_64_) );
	NOR2X1 NOR2X1_200 ( .A(target[2]), .B(Y_10_), .Y(_65_) );
	OAI22X1 OAI22X1_213 ( .A(_61_), .B(_62_), .C(_64_), .D(_65_), .Y(_66_) );
	INVX1 INVX1_311 ( .A(Y_11_), .Y(_67_) );
	NOR2X1 NOR2X1_201 ( .A(target[3]), .B(_67_), .Y(_68_) );
	NAND2X1 NAND2X1_318 ( .A(target[3]), .B(_67_), .Y(_69_) );
	INVX1 INVX1_312 ( .A(Y_10_), .Y(_70_) );
	NOR2X1 NOR2X1_202 ( .A(target[2]), .B(_70_), .Y(_71_) );
	AOI21X1 AOI21X1_254 ( .A(_69_), .B(_71_), .C(_68_), .Y(_72_) );
	OAI21X1 OAI21X1_401 ( .A(_66_), .B(_59_), .C(_72_), .Y(_73_) );
	INVX1 INVX1_313 ( .A(Y_14_), .Y(_74_) );
	NAND2X1 NAND2X1_319 ( .A(target[6]), .B(_74_), .Y(_75_) );
	INVX1 INVX1_314 ( .A(Y_15_), .Y(_76_) );
	NAND2X1 NAND2X1_320 ( .A(target[7]), .B(_76_), .Y(_77_) );
	INVX1 INVX1_315 ( .A(target[6]), .Y(_78_) );
	AOI22X1 AOI22X1_6 ( .A(_45_), .B(Y_15_), .C(_78_), .D(Y_14_), .Y(_79_) );
	NAND3X1 NAND3X1_63 ( .A(_75_), .B(_77_), .C(_79_), .Y(_80_) );
	AOI22X1 AOI22X1_7 ( .A(_37_), .B(Y_13_), .C(_38_), .D(Y_12_), .Y(_81_) );
	INVX1 INVX1_316 ( .A(Y_13_), .Y(_82_) );
	INVX1 INVX1_317 ( .A(Y_12_), .Y(_83_) );
	AOI22X1 AOI22X1_8 ( .A(_82_), .B(target[5]), .C(target[4]), .D(_83_), .Y(_84_) );
	NAND2X1 NAND2X1_321 ( .A(_81_), .B(_84_), .Y(_85_) );
	NOR2X1 NOR2X1_203 ( .A(_85_), .B(_80_), .Y(_86_) );
	OAI22X1 OAI22X1_214 ( .A(_82_), .B(target[5]), .C(target[4]), .D(_83_), .Y(_87_) );
	OAI21X1 OAI21X1_402 ( .A(_37_), .B(Y_13_), .C(_87_), .Y(_88_) );
	OAI22X1 OAI22X1_215 ( .A(_76_), .B(target[7]), .C(target[6]), .D(_74_), .Y(_89_) );
	AOI21X1 AOI21X1_255 ( .A(_77_), .B(_89_), .C(_1__bF_buf1), .Y(_90_) );
	OAI21X1 OAI21X1_403 ( .A(_80_), .B(_88_), .C(_90_), .Y(_91_) );
	AOI21X1 AOI21X1_256 ( .A(_73_), .B(_86_), .C(_91_), .Y(_92_) );
	NAND3X1 NAND3X1_64 ( .A(Y_0_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_93_) );
	INVX1 INVX1_318 ( .A(target[1]), .Y(_94_) );
	NAND2X1 NAND2X1_322 ( .A(Y_17_), .B(_94_), .Y(_95_) );
	INVX1 INVX1_319 ( .A(target[0]), .Y(_96_) );
	OAI22X1 OAI22X1_216 ( .A(_94_), .B(Y_17_), .C(_96_), .D(Y_16_), .Y(_97_) );
	NAND2X1 NAND2X1_323 ( .A(_95_), .B(_97_), .Y(_98_) );
	NAND2X1 NAND2X1_324 ( .A(target[3]), .B(Y_19_), .Y(_99_) );
	OR2X2 OR2X2_19 ( .A(target[3]), .B(Y_19_), .Y(_100_) );
	INVX1 INVX1_320 ( .A(target[2]), .Y(_101_) );
	NAND2X1 NAND2X1_325 ( .A(_101_), .B(_26_), .Y(_102_) );
	AOI22X1 AOI22X1_9 ( .A(_99_), .B(_100_), .C(_102_), .D(_19_), .Y(_103_) );
	INVX1 INVX1_321 ( .A(target[3]), .Y(_104_) );
	NAND2X1 NAND2X1_326 ( .A(Y_19_), .B(_104_), .Y(_105_) );
	NOR2X1 NOR2X1_204 ( .A(Y_19_), .B(_104_), .Y(_106_) );
	NAND2X1 NAND2X1_327 ( .A(Y_18_), .B(_101_), .Y(_107_) );
	OAI21X1 OAI21X1_404 ( .A(_106_), .B(_107_), .C(_105_), .Y(_108_) );
	AOI21X1 AOI21X1_257 ( .A(_103_), .B(_98_), .C(_108_), .Y(_109_) );
	NAND2X1 NAND2X1_328 ( .A(_45_), .B(_46_), .Y(_110_) );
	NAND2X1 NAND2X1_329 ( .A(_78_), .B(_47_), .Y(_111_) );
	AOI22X1 AOI22X1_10 ( .A(_110_), .B(_30_), .C(_33_), .D(_111_), .Y(_112_) );
	NAND3X1 NAND3X1_65 ( .A(_39_), .B(_42_), .C(_112_), .Y(_113_) );
	NAND2X1 NAND2X1_330 ( .A(target[7]), .B(_46_), .Y(_114_) );
	AOI21X1 AOI21X1_258 ( .A(target[5]), .B(_40_), .C(_39_), .Y(_115_) );
	AOI22X1 AOI22X1_11 ( .A(_114_), .B(_48_), .C(_115_), .D(_112_), .Y(_116_) );
	OAI21X1 OAI21X1_405 ( .A(_109_), .B(_113_), .C(_116_), .Y(_117_) );
	NAND2X1 NAND2X1_331 ( .A(Y_9_), .B(_94_), .Y(_118_) );
	OAI22X1 OAI22X1_217 ( .A(_94_), .B(Y_9_), .C(Y_8_), .D(_96_), .Y(_119_) );
	NAND2X1 NAND2X1_332 ( .A(_118_), .B(_119_), .Y(_120_) );
	OR2X2 OR2X2_20 ( .A(target[3]), .B(Y_11_), .Y(_121_) );
	NAND2X1 NAND2X1_333 ( .A(_101_), .B(_70_), .Y(_122_) );
	AOI22X1 AOI22X1_12 ( .A(_60_), .B(_121_), .C(_122_), .D(_63_), .Y(_123_) );
	NAND2X1 NAND2X1_334 ( .A(Y_11_), .B(_104_), .Y(_124_) );
	NOR2X1 NOR2X1_205 ( .A(Y_11_), .B(_104_), .Y(_125_) );
	NAND2X1 NAND2X1_335 ( .A(Y_10_), .B(_101_), .Y(_126_) );
	OAI21X1 OAI21X1_406 ( .A(_125_), .B(_126_), .C(_124_), .Y(_127_) );
	AOI21X1 AOI21X1_259 ( .A(_123_), .B(_120_), .C(_127_), .Y(_128_) );
	NAND2X1 NAND2X1_336 ( .A(target[6]), .B(Y_14_), .Y(_129_) );
	NAND2X1 NAND2X1_337 ( .A(_78_), .B(_74_), .Y(_130_) );
	NAND2X1 NAND2X1_338 ( .A(target[7]), .B(Y_15_), .Y(_131_) );
	NAND2X1 NAND2X1_339 ( .A(_45_), .B(_76_), .Y(_132_) );
	AOI22X1 AOI22X1_13 ( .A(_130_), .B(_129_), .C(_131_), .D(_132_), .Y(_133_) );
	OAI22X1 OAI22X1_218 ( .A(_37_), .B(Y_13_), .C(_38_), .D(Y_12_), .Y(_134_) );
	NOR2X1 NOR2X1_206 ( .A(_87_), .B(_134_), .Y(_135_) );
	NAND2X1 NAND2X1_340 ( .A(_133_), .B(_135_), .Y(_136_) );
	AOI21X1 AOI21X1_260 ( .A(target[5]), .B(_82_), .C(_81_), .Y(_137_) );
	INVX1 INVX1_322 ( .A(_1__bF_buf0), .Y(_138_) );
	NOR2X1 NOR2X1_207 ( .A(Y_15_), .B(_45_), .Y(_139_) );
	OAI21X1 OAI21X1_407 ( .A(_79_), .B(_139_), .C(_138_), .Y(_140_) );
	AOI21X1 AOI21X1_261 ( .A(_133_), .B(_137_), .C(_140_), .Y(_141_) );
	OAI21X1 OAI21X1_408 ( .A(_128_), .B(_136_), .C(_141_), .Y(_142_) );
	OAI21X1 OAI21X1_409 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(bounty_synth_0_), .Y(_143_) );
	AOI21X1 AOI21X1_262 ( .A(_93_), .B(_143_), .C(_10__bF_buf6), .Y(_7__0_) );
	NAND3X1 NAND3X1_66 ( .A(Y_1_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_144_) );
	OAI21X1 OAI21X1_410 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(bounty_synth_1_), .Y(_145_) );
	AOI21X1 AOI21X1_263 ( .A(_144_), .B(_145_), .C(_10__bF_buf5), .Y(_7__1_) );
	NAND3X1 NAND3X1_67 ( .A(Y_2_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_146_) );
	OAI21X1 OAI21X1_411 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(bounty_synth_2_), .Y(_147_) );
	AOI21X1 AOI21X1_264 ( .A(_146_), .B(_147_), .C(_10__bF_buf4), .Y(_7__2_) );
	NAND3X1 NAND3X1_68 ( .A(Y_3_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_148_) );
	OAI21X1 OAI21X1_412 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(bounty_synth_3_), .Y(_149_) );
	AOI21X1 AOI21X1_265 ( .A(_148_), .B(_149_), .C(_10__bF_buf3), .Y(_7__3_) );
	NAND3X1 NAND3X1_69 ( .A(Y_4_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_150_) );
	OAI21X1 OAI21X1_413 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(bounty_synth_4_), .Y(_151_) );
	AOI21X1 AOI21X1_266 ( .A(_150_), .B(_151_), .C(_10__bF_buf2), .Y(_7__4_) );
	NAND3X1 NAND3X1_70 ( .A(Y_5_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_152_) );
	OAI21X1 OAI21X1_414 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(bounty_synth_5_), .Y(_153_) );
	AOI21X1 AOI21X1_267 ( .A(_152_), .B(_153_), .C(_10__bF_buf1), .Y(_7__5_) );
	NAND3X1 NAND3X1_71 ( .A(Y_6_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_154_) );
	OAI21X1 OAI21X1_415 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(bounty_synth_6_), .Y(_155_) );
	AOI21X1 AOI21X1_268 ( .A(_154_), .B(_155_), .C(_10__bF_buf0), .Y(_7__6_) );
	NAND3X1 NAND3X1_72 ( .A(Y_7_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_156_) );
	OAI21X1 OAI21X1_416 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(bounty_synth_7_), .Y(_157_) );
	AOI21X1 AOI21X1_269 ( .A(_156_), .B(_157_), .C(_10__bF_buf6), .Y(_7__7_) );
	NAND3X1 NAND3X1_73 ( .A(Y_8_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_158_) );
	OAI21X1 OAI21X1_417 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(bounty_synth_8_), .Y(_159_) );
	AOI21X1 AOI21X1_270 ( .A(_158_), .B(_159_), .C(_10__bF_buf5), .Y(_7__8_) );
	NAND3X1 NAND3X1_74 ( .A(Y_9_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_160_) );
	OAI21X1 OAI21X1_418 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(bounty_synth_9_), .Y(_161_) );
	AOI21X1 AOI21X1_271 ( .A(_160_), .B(_161_), .C(_10__bF_buf4), .Y(_7__9_) );
	NAND3X1 NAND3X1_75 ( .A(Y_10_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_162_) );
	OAI21X1 OAI21X1_419 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(bounty_synth_10_), .Y(_163_) );
	AOI21X1 AOI21X1_272 ( .A(_162_), .B(_163_), .C(_10__bF_buf3), .Y(_7__10_) );
	NAND3X1 NAND3X1_76 ( .A(Y_11_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_164_) );
	OAI21X1 OAI21X1_420 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(bounty_synth_11_), .Y(_165_) );
	AOI21X1 AOI21X1_273 ( .A(_164_), .B(_165_), .C(_10__bF_buf2), .Y(_7__11_) );
	NAND3X1 NAND3X1_77 ( .A(Y_12_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_166_) );
	OAI21X1 OAI21X1_421 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(bounty_synth_12_), .Y(_167_) );
	AOI21X1 AOI21X1_274 ( .A(_166_), .B(_167_), .C(_10__bF_buf1), .Y(_7__12_) );
	NAND3X1 NAND3X1_78 ( .A(Y_13_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_168_) );
	OAI21X1 OAI21X1_422 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(bounty_synth_13_), .Y(_169_) );
	AOI21X1 AOI21X1_275 ( .A(_168_), .B(_169_), .C(_10__bF_buf0), .Y(_7__13_) );
	NAND3X1 NAND3X1_79 ( .A(Y_14_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_170_) );
	OAI21X1 OAI21X1_423 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(bounty_synth_14_), .Y(_171_) );
	AOI21X1 AOI21X1_276 ( .A(_170_), .B(_171_), .C(_10__bF_buf6), .Y(_7__14_) );
	NAND3X1 NAND3X1_80 ( .A(Y_15_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_172_) );
	OAI21X1 OAI21X1_424 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(bounty_synth_15_), .Y(_173_) );
	AOI21X1 AOI21X1_277 ( .A(_172_), .B(_173_), .C(_10__bF_buf5), .Y(_7__15_) );
	NAND3X1 NAND3X1_81 ( .A(Y_16_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_174_) );
	OAI21X1 OAI21X1_425 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(bounty_synth_16_), .Y(_175_) );
	AOI21X1 AOI21X1_278 ( .A(_174_), .B(_175_), .C(_10__bF_buf4), .Y(_7__16_) );
	NAND3X1 NAND3X1_82 ( .A(Y_17_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_176_) );
	OAI21X1 OAI21X1_426 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(bounty_synth_17_), .Y(_177_) );
	AOI21X1 AOI21X1_279 ( .A(_176_), .B(_177_), .C(_10__bF_buf3), .Y(_7__17_) );
	NAND3X1 NAND3X1_83 ( .A(Y_18_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_178_) );
	OAI21X1 OAI21X1_427 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(bounty_synth_18_), .Y(_179_) );
	AOI21X1 AOI21X1_280 ( .A(_178_), .B(_179_), .C(_10__bF_buf2), .Y(_7__18_) );
	NAND3X1 NAND3X1_84 ( .A(Y_19_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_180_) );
	OAI21X1 OAI21X1_428 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(bounty_synth_19_), .Y(_181_) );
	AOI21X1 AOI21X1_281 ( .A(_180_), .B(_181_), .C(_10__bF_buf1), .Y(_7__19_) );
	NAND3X1 NAND3X1_85 ( .A(Y_20_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_182_) );
	OAI21X1 OAI21X1_429 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(bounty_synth_20_), .Y(_183_) );
	AOI21X1 AOI21X1_282 ( .A(_182_), .B(_183_), .C(_10__bF_buf0), .Y(_7__20_) );
	NAND3X1 NAND3X1_86 ( .A(Y_21_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_184_) );
	OAI21X1 OAI21X1_430 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(bounty_synth_21_), .Y(_185_) );
	AOI21X1 AOI21X1_283 ( .A(_184_), .B(_185_), .C(_10__bF_buf6), .Y(_7__21_) );
	NAND3X1 NAND3X1_87 ( .A(Y_22_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_186_) );
	OAI21X1 OAI21X1_431 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(bounty_synth_22_), .Y(_187_) );
	AOI21X1 AOI21X1_284 ( .A(_186_), .B(_187_), .C(_10__bF_buf5), .Y(_7__22_) );
	NAND3X1 NAND3X1_88 ( .A(Y_23_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_188_) );
	OAI21X1 OAI21X1_432 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(bounty_synth_23_), .Y(_189_) );
	AOI21X1 AOI21X1_285 ( .A(_188_), .B(_189_), .C(_10__bF_buf4), .Y(_7__23_) );
	NAND3X1 NAND3X1_89 ( .A(Ynonce_synth_0_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_190_) );
	OAI21X1 OAI21X1_433 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_0_), .Y(_191_) );
	AOI21X1 AOI21X1_286 ( .A(_190_), .B(_191_), .C(_10__bF_buf3), .Y(_8__0_) );
	NAND3X1 NAND3X1_90 ( .A(Ynonce_synth_1_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_192_) );
	OAI21X1 OAI21X1_434 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_1_), .Y(_193_) );
	AOI21X1 AOI21X1_287 ( .A(_192_), .B(_193_), .C(_10__bF_buf2), .Y(_8__1_) );
	NAND3X1 NAND3X1_91 ( .A(Ynonce_synth_2_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_194_) );
	OAI21X1 OAI21X1_435 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_2_), .Y(_195_) );
	AOI21X1 AOI21X1_288 ( .A(_194_), .B(_195_), .C(_10__bF_buf1), .Y(_8__2_) );
	NAND3X1 NAND3X1_92 ( .A(Ynonce_synth_3_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_196_) );
	OAI21X1 OAI21X1_436 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_3_), .Y(_197_) );
	AOI21X1 AOI21X1_289 ( .A(_196_), .B(_197_), .C(_10__bF_buf0), .Y(_8__3_) );
	NAND3X1 NAND3X1_93 ( .A(Ynonce_synth_4_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_198_) );
	OAI21X1 OAI21X1_437 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(comparador_nonce_synth_valido_4_), .Y(_199_) );
	AOI21X1 AOI21X1_290 ( .A(_198_), .B(_199_), .C(_10__bF_buf6), .Y(_8__4_) );
	NAND3X1 NAND3X1_94 ( .A(Ynonce_synth_5_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_200_) );
	OAI21X1 OAI21X1_438 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(comparador_nonce_synth_valido_5_), .Y(_201_) );
	AOI21X1 AOI21X1_291 ( .A(_200_), .B(_201_), .C(_10__bF_buf5), .Y(_8__5_) );
	NAND3X1 NAND3X1_95 ( .A(Ynonce_synth_6_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_202_) );
	OAI21X1 OAI21X1_439 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(comparador_nonce_synth_valido_6_), .Y(_203_) );
	AOI21X1 AOI21X1_292 ( .A(_202_), .B(_203_), .C(_10__bF_buf4), .Y(_8__6_) );
	NAND3X1 NAND3X1_96 ( .A(Ynonce_synth_7_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_204_) );
	OAI21X1 OAI21X1_440 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_7_), .Y(_205_) );
	AOI21X1 AOI21X1_293 ( .A(_204_), .B(_205_), .C(_10__bF_buf3), .Y(_8__7_) );
	NAND3X1 NAND3X1_97 ( .A(Ynonce_synth_8_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_206_) );
	OAI21X1 OAI21X1_441 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_8_), .Y(_207_) );
	AOI21X1 AOI21X1_294 ( .A(_206_), .B(_207_), .C(_10__bF_buf2), .Y(_8__8_) );
	NAND3X1 NAND3X1_98 ( .A(Ynonce_synth_9_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_208_) );
	OAI21X1 OAI21X1_442 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_9_), .Y(_209_) );
	AOI21X1 AOI21X1_295 ( .A(_208_), .B(_209_), .C(_10__bF_buf1), .Y(_8__9_) );
	NAND3X1 NAND3X1_99 ( .A(Ynonce_synth_10_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_210_) );
	OAI21X1 OAI21X1_443 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_10_), .Y(_211_) );
	AOI21X1 AOI21X1_296 ( .A(_210_), .B(_211_), .C(_10__bF_buf0), .Y(_8__10_) );
	NAND3X1 NAND3X1_100 ( .A(Ynonce_synth_11_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_212_) );
	OAI21X1 OAI21X1_444 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(comparador_nonce_synth_valido_11_), .Y(_213_) );
	AOI21X1 AOI21X1_297 ( .A(_212_), .B(_213_), .C(_10__bF_buf6), .Y(_8__11_) );
	NAND3X1 NAND3X1_101 ( .A(Ynonce_synth_12_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_214_) );
	OAI21X1 OAI21X1_445 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(comparador_nonce_synth_valido_12_), .Y(_215_) );
	AOI21X1 AOI21X1_298 ( .A(_214_), .B(_215_), .C(_10__bF_buf5), .Y(_8__12_) );
	NAND3X1 NAND3X1_102 ( .A(Ynonce_synth_13_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_216_) );
	OAI21X1 OAI21X1_446 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(comparador_nonce_synth_valido_13_), .Y(_217_) );
	AOI21X1 AOI21X1_299 ( .A(_216_), .B(_217_), .C(_10__bF_buf4), .Y(_8__13_) );
	NAND3X1 NAND3X1_103 ( .A(Ynonce_synth_14_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_218_) );
	OAI21X1 OAI21X1_447 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_14_), .Y(_219_) );
	AOI21X1 AOI21X1_300 ( .A(_218_), .B(_219_), .C(_10__bF_buf3), .Y(_8__14_) );
	NAND3X1 NAND3X1_104 ( .A(Ynonce_synth_15_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_220_) );
	OAI21X1 OAI21X1_448 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_15_), .Y(_221_) );
	AOI21X1 AOI21X1_301 ( .A(_220_), .B(_221_), .C(_10__bF_buf2), .Y(_8__15_) );
	NAND3X1 NAND3X1_105 ( .A(Ynonce_synth_16_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_222_) );
	OAI21X1 OAI21X1_449 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_16_), .Y(_223_) );
	AOI21X1 AOI21X1_302 ( .A(_222_), .B(_223_), .C(_10__bF_buf1), .Y(_8__16_) );
	NAND3X1 NAND3X1_106 ( .A(Ynonce_synth_17_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_224_) );
	OAI21X1 OAI21X1_450 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_17_), .Y(_225_) );
	AOI21X1 AOI21X1_303 ( .A(_224_), .B(_225_), .C(_10__bF_buf0), .Y(_8__17_) );
	NAND3X1 NAND3X1_107 ( .A(Ynonce_synth_18_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_226_) );
	OAI21X1 OAI21X1_451 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(comparador_nonce_synth_valido_18_), .Y(_227_) );
	AOI21X1 AOI21X1_304 ( .A(_226_), .B(_227_), .C(_10__bF_buf6), .Y(_8__18_) );
	NAND3X1 NAND3X1_108 ( .A(Ynonce_synth_19_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_228_) );
	OAI21X1 OAI21X1_452 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(comparador_nonce_synth_valido_19_), .Y(_229_) );
	AOI21X1 AOI21X1_305 ( .A(_228_), .B(_229_), .C(_10__bF_buf5), .Y(_8__19_) );
	NAND3X1 NAND3X1_109 ( .A(Ynonce_synth_20_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_230_) );
	OAI21X1 OAI21X1_453 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(comparador_nonce_synth_valido_20_), .Y(_231_) );
	AOI21X1 AOI21X1_306 ( .A(_230_), .B(_231_), .C(_10__bF_buf4), .Y(_8__20_) );
	NAND3X1 NAND3X1_110 ( .A(Ynonce_synth_21_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_232_) );
	OAI21X1 OAI21X1_454 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_21_), .Y(_233_) );
	AOI21X1 AOI21X1_307 ( .A(_232_), .B(_233_), .C(_10__bF_buf3), .Y(_8__21_) );
	NAND3X1 NAND3X1_111 ( .A(Ynonce_synth_22_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_234_) );
	OAI21X1 OAI21X1_455 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_22_), .Y(_235_) );
	AOI21X1 AOI21X1_308 ( .A(_234_), .B(_235_), .C(_10__bF_buf2), .Y(_8__22_) );
	NAND3X1 NAND3X1_112 ( .A(Ynonce_synth_23_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_236_) );
	OAI21X1 OAI21X1_456 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_23_), .Y(_237_) );
	AOI21X1 AOI21X1_309 ( .A(_236_), .B(_237_), .C(_10__bF_buf1), .Y(_8__23_) );
	NAND3X1 NAND3X1_113 ( .A(Ynonce_synth_24_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_238_) );
	OAI21X1 OAI21X1_457 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_24_), .Y(_239_) );
	AOI21X1 AOI21X1_310 ( .A(_238_), .B(_239_), .C(_10__bF_buf0), .Y(_8__24_) );
	NAND3X1 NAND3X1_114 ( .A(Ynonce_synth_25_), .B(_53__bF_buf6), .C(_92__bF_buf6), .Y(_240_) );
	OAI21X1 OAI21X1_458 ( .A(_117__bF_buf6), .B(_142__bF_buf6), .C(comparador_nonce_synth_valido_25_), .Y(_241_) );
	AOI21X1 AOI21X1_311 ( .A(_240_), .B(_241_), .C(_10__bF_buf6), .Y(_8__25_) );
	NAND3X1 NAND3X1_115 ( .A(Ynonce_synth_26_), .B(_53__bF_buf5), .C(_92__bF_buf5), .Y(_242_) );
	OAI21X1 OAI21X1_459 ( .A(_117__bF_buf5), .B(_142__bF_buf5), .C(comparador_nonce_synth_valido_26_), .Y(_243_) );
	AOI21X1 AOI21X1_312 ( .A(_242_), .B(_243_), .C(_10__bF_buf5), .Y(_8__26_) );
	NAND3X1 NAND3X1_116 ( .A(Ynonce_synth_27_), .B(_53__bF_buf4), .C(_92__bF_buf4), .Y(_244_) );
	OAI21X1 OAI21X1_460 ( .A(_117__bF_buf4), .B(_142__bF_buf4), .C(comparador_nonce_synth_valido_27_), .Y(_245_) );
	AOI21X1 AOI21X1_313 ( .A(_244_), .B(_245_), .C(_10__bF_buf4), .Y(_8__27_) );
	NAND3X1 NAND3X1_117 ( .A(Ynonce_synth_28_), .B(_53__bF_buf3), .C(_92__bF_buf3), .Y(_246_) );
	OAI21X1 OAI21X1_461 ( .A(_117__bF_buf3), .B(_142__bF_buf3), .C(comparador_nonce_synth_valido_28_), .Y(_247_) );
	AOI21X1 AOI21X1_314 ( .A(_246_), .B(_247_), .C(_10__bF_buf3), .Y(_8__28_) );
	NAND3X1 NAND3X1_118 ( .A(Ynonce_synth_29_), .B(_53__bF_buf2), .C(_92__bF_buf2), .Y(_248_) );
	OAI21X1 OAI21X1_462 ( .A(_117__bF_buf2), .B(_142__bF_buf2), .C(comparador_nonce_synth_valido_29_), .Y(_249_) );
	AOI21X1 AOI21X1_315 ( .A(_248_), .B(_249_), .C(_10__bF_buf2), .Y(_8__29_) );
	NAND3X1 NAND3X1_119 ( .A(Ynonce_synth_30_), .B(_53__bF_buf1), .C(_92__bF_buf1), .Y(_250_) );
	OAI21X1 OAI21X1_463 ( .A(_117__bF_buf1), .B(_142__bF_buf1), .C(comparador_nonce_synth_valido_30_), .Y(_251_) );
	AOI21X1 AOI21X1_316 ( .A(_250_), .B(_251_), .C(_10__bF_buf1), .Y(_8__30_) );
	NAND3X1 NAND3X1_120 ( .A(Ynonce_synth_31_), .B(_53__bF_buf0), .C(_92__bF_buf0), .Y(_252_) );
	OAI21X1 OAI21X1_464 ( .A(_117__bF_buf0), .B(_142__bF_buf0), .C(comparador_nonce_synth_valido_31_), .Y(_253_) );
	AOI21X1 AOI21X1_317 ( .A(_252_), .B(_253_), .C(_10__bF_buf0), .Y(_8__31_) );
	AOI21X1 AOI21X1_318 ( .A(_53__bF_buf6), .B(_92__bF_buf6), .C(comparador_valid_bF_buf2), .Y(_254_) );
	OAI21X1 OAI21X1_465 ( .A(_53__bF_buf5), .B(_1__bF_buf5), .C(reset_L_bF_buf43), .Y(_255_) );
	NOR2X1 NOR2X1_208 ( .A(_255_), .B(_254_), .Y(_9_) );
	DFFPOSX1 DFFPOSX1_484 ( .CLK(clk_bF_buf86), .D(_9_), .Q(comparador_valid) );
	DFFPOSX1 DFFPOSX1_485 ( .CLK(clk_bF_buf85), .D(_8__0_), .Q(comparador_nonce_synth_valido_0_) );
	DFFPOSX1 DFFPOSX1_486 ( .CLK(clk_bF_buf84), .D(_8__1_), .Q(comparador_nonce_synth_valido_1_) );
	DFFPOSX1 DFFPOSX1_487 ( .CLK(clk_bF_buf83), .D(_8__2_), .Q(comparador_nonce_synth_valido_2_) );
	DFFPOSX1 DFFPOSX1_488 ( .CLK(clk_bF_buf82), .D(_8__3_), .Q(comparador_nonce_synth_valido_3_) );
	DFFPOSX1 DFFPOSX1_489 ( .CLK(clk_bF_buf81), .D(_8__4_), .Q(comparador_nonce_synth_valido_4_) );
	DFFPOSX1 DFFPOSX1_490 ( .CLK(clk_bF_buf80), .D(_8__5_), .Q(comparador_nonce_synth_valido_5_) );
	DFFPOSX1 DFFPOSX1_491 ( .CLK(clk_bF_buf79), .D(_8__6_), .Q(comparador_nonce_synth_valido_6_) );
	DFFPOSX1 DFFPOSX1_492 ( .CLK(clk_bF_buf78), .D(_8__7_), .Q(comparador_nonce_synth_valido_7_) );
	DFFPOSX1 DFFPOSX1_493 ( .CLK(clk_bF_buf77), .D(_8__8_), .Q(comparador_nonce_synth_valido_8_) );
	DFFPOSX1 DFFPOSX1_494 ( .CLK(clk_bF_buf76), .D(_8__9_), .Q(comparador_nonce_synth_valido_9_) );
	DFFPOSX1 DFFPOSX1_495 ( .CLK(clk_bF_buf75), .D(_8__10_), .Q(comparador_nonce_synth_valido_10_) );
	DFFPOSX1 DFFPOSX1_496 ( .CLK(clk_bF_buf74), .D(_8__11_), .Q(comparador_nonce_synth_valido_11_) );
	DFFPOSX1 DFFPOSX1_497 ( .CLK(clk_bF_buf73), .D(_8__12_), .Q(comparador_nonce_synth_valido_12_) );
	DFFPOSX1 DFFPOSX1_498 ( .CLK(clk_bF_buf72), .D(_8__13_), .Q(comparador_nonce_synth_valido_13_) );
	DFFPOSX1 DFFPOSX1_499 ( .CLK(clk_bF_buf71), .D(_8__14_), .Q(comparador_nonce_synth_valido_14_) );
	DFFPOSX1 DFFPOSX1_500 ( .CLK(clk_bF_buf70), .D(_8__15_), .Q(comparador_nonce_synth_valido_15_) );
	DFFPOSX1 DFFPOSX1_501 ( .CLK(clk_bF_buf69), .D(_8__16_), .Q(comparador_nonce_synth_valido_16_) );
	DFFPOSX1 DFFPOSX1_502 ( .CLK(clk_bF_buf68), .D(_8__17_), .Q(comparador_nonce_synth_valido_17_) );
	DFFPOSX1 DFFPOSX1_503 ( .CLK(clk_bF_buf67), .D(_8__18_), .Q(comparador_nonce_synth_valido_18_) );
	DFFPOSX1 DFFPOSX1_504 ( .CLK(clk_bF_buf66), .D(_8__19_), .Q(comparador_nonce_synth_valido_19_) );
	DFFPOSX1 DFFPOSX1_505 ( .CLK(clk_bF_buf65), .D(_8__20_), .Q(comparador_nonce_synth_valido_20_) );
	DFFPOSX1 DFFPOSX1_506 ( .CLK(clk_bF_buf64), .D(_8__21_), .Q(comparador_nonce_synth_valido_21_) );
	DFFPOSX1 DFFPOSX1_507 ( .CLK(clk_bF_buf63), .D(_8__22_), .Q(comparador_nonce_synth_valido_22_) );
	DFFPOSX1 DFFPOSX1_508 ( .CLK(clk_bF_buf62), .D(_8__23_), .Q(comparador_nonce_synth_valido_23_) );
	DFFPOSX1 DFFPOSX1_509 ( .CLK(clk_bF_buf61), .D(_8__24_), .Q(comparador_nonce_synth_valido_24_) );
	DFFPOSX1 DFFPOSX1_510 ( .CLK(clk_bF_buf60), .D(_8__25_), .Q(comparador_nonce_synth_valido_25_) );
	DFFPOSX1 DFFPOSX1_511 ( .CLK(clk_bF_buf59), .D(_8__26_), .Q(comparador_nonce_synth_valido_26_) );
	DFFPOSX1 DFFPOSX1_512 ( .CLK(clk_bF_buf58), .D(_8__27_), .Q(comparador_nonce_synth_valido_27_) );
	DFFPOSX1 DFFPOSX1_513 ( .CLK(clk_bF_buf57), .D(_8__28_), .Q(comparador_nonce_synth_valido_28_) );
	DFFPOSX1 DFFPOSX1_514 ( .CLK(clk_bF_buf56), .D(_8__29_), .Q(comparador_nonce_synth_valido_29_) );
	DFFPOSX1 DFFPOSX1_515 ( .CLK(clk_bF_buf55), .D(_8__30_), .Q(comparador_nonce_synth_valido_30_) );
	DFFPOSX1 DFFPOSX1_516 ( .CLK(clk_bF_buf54), .D(_8__31_), .Q(comparador_nonce_synth_valido_31_) );
	DFFPOSX1 DFFPOSX1_517 ( .CLK(clk_bF_buf53), .D(_7__0_), .Q(bounty_synth_0_) );
	DFFPOSX1 DFFPOSX1_518 ( .CLK(clk_bF_buf52), .D(_7__1_), .Q(bounty_synth_1_) );
	DFFPOSX1 DFFPOSX1_519 ( .CLK(clk_bF_buf51), .D(_7__2_), .Q(bounty_synth_2_) );
	DFFPOSX1 DFFPOSX1_520 ( .CLK(clk_bF_buf50), .D(_7__3_), .Q(bounty_synth_3_) );
	DFFPOSX1 DFFPOSX1_521 ( .CLK(clk_bF_buf49), .D(_7__4_), .Q(bounty_synth_4_) );
	DFFPOSX1 DFFPOSX1_522 ( .CLK(clk_bF_buf48), .D(_7__5_), .Q(bounty_synth_5_) );
	DFFPOSX1 DFFPOSX1_523 ( .CLK(clk_bF_buf47), .D(_7__6_), .Q(bounty_synth_6_) );
	DFFPOSX1 DFFPOSX1_524 ( .CLK(clk_bF_buf46), .D(_7__7_), .Q(bounty_synth_7_) );
	DFFPOSX1 DFFPOSX1_525 ( .CLK(clk_bF_buf45), .D(_7__8_), .Q(bounty_synth_8_) );
	DFFPOSX1 DFFPOSX1_526 ( .CLK(clk_bF_buf44), .D(_7__9_), .Q(bounty_synth_9_) );
	DFFPOSX1 DFFPOSX1_527 ( .CLK(clk_bF_buf43), .D(_7__10_), .Q(bounty_synth_10_) );
	DFFPOSX1 DFFPOSX1_528 ( .CLK(clk_bF_buf42), .D(_7__11_), .Q(bounty_synth_11_) );
	DFFPOSX1 DFFPOSX1_529 ( .CLK(clk_bF_buf41), .D(_7__12_), .Q(bounty_synth_12_) );
	DFFPOSX1 DFFPOSX1_530 ( .CLK(clk_bF_buf40), .D(_7__13_), .Q(bounty_synth_13_) );
	DFFPOSX1 DFFPOSX1_531 ( .CLK(clk_bF_buf39), .D(_7__14_), .Q(bounty_synth_14_) );
	DFFPOSX1 DFFPOSX1_532 ( .CLK(clk_bF_buf38), .D(_7__15_), .Q(bounty_synth_15_) );
	DFFPOSX1 DFFPOSX1_533 ( .CLK(clk_bF_buf37), .D(_7__16_), .Q(bounty_synth_16_) );
	DFFPOSX1 DFFPOSX1_534 ( .CLK(clk_bF_buf36), .D(_7__17_), .Q(bounty_synth_17_) );
	DFFPOSX1 DFFPOSX1_535 ( .CLK(clk_bF_buf35), .D(_7__18_), .Q(bounty_synth_18_) );
	DFFPOSX1 DFFPOSX1_536 ( .CLK(clk_bF_buf34), .D(_7__19_), .Q(bounty_synth_19_) );
	DFFPOSX1 DFFPOSX1_537 ( .CLK(clk_bF_buf33), .D(_7__20_), .Q(bounty_synth_20_) );
	DFFPOSX1 DFFPOSX1_538 ( .CLK(clk_bF_buf32), .D(_7__21_), .Q(bounty_synth_21_) );
	DFFPOSX1 DFFPOSX1_539 ( .CLK(clk_bF_buf31), .D(_7__22_), .Q(bounty_synth_22_) );
	DFFPOSX1 DFFPOSX1_540 ( .CLK(clk_bF_buf30), .D(_7__23_), .Q(bounty_synth_23_) );
	INVX1 INVX1_323 ( .A(bloque_in_1_32_), .Y(_546_) );
	NOR2X1 NOR2X1_209 ( .A(concatenador_counter_2d_1_bF_buf0), .B(concatenador_counter_2d_0_bF_buf8), .Y(_547_) );
	NOR2X1 NOR2X1_210 ( .A(concatenador_counter_2d_3_), .B(concatenador_counter_2d_2_), .Y(_548_) );
	NOR2X1 NOR2X1_211 ( .A(concatenador_counter_2d_5_), .B(concatenador_counter_2d_4_), .Y(_549_) );
	NAND3X1 NAND3X1_121 ( .A(_547_), .B(_548_), .C(_549_), .Y(_550_) );
	OAI21X1 OAI21X1_466 ( .A(_550__bF_buf15), .B(RAM_entrada_89_), .C(reset_L_bF_buf42), .Y(_551_) );
	AOI21X1 AOI21X1_319 ( .A(_546_), .B(_550__bF_buf14), .C(_551_), .Y(_257__32_) );
	INVX1 INVX1_324 ( .A(bloque_in_1_33_), .Y(_552_) );
	OAI21X1 OAI21X1_467 ( .A(_550__bF_buf13), .B(RAM_entrada_77_), .C(reset_L_bF_buf41), .Y(_553_) );
	AOI21X1 AOI21X1_320 ( .A(_552_), .B(_550__bF_buf12), .C(_553_), .Y(_257__33_) );
	INVX1 INVX1_325 ( .A(bloque_in_1_34_), .Y(_554_) );
	OAI21X1 OAI21X1_468 ( .A(_550__bF_buf11), .B(RAM_entrada_84_bF_buf3), .C(reset_L_bF_buf40), .Y(_555_) );
	AOI21X1 AOI21X1_321 ( .A(_554_), .B(_550__bF_buf10), .C(_555_), .Y(_257__34_) );
	INVX1 INVX1_326 ( .A(bloque_in_1_35_), .Y(_556_) );
	OAI21X1 OAI21X1_469 ( .A(_550__bF_buf9), .B(RAM_entrada_94_), .C(reset_L_bF_buf39), .Y(_557_) );
	AOI21X1 AOI21X1_322 ( .A(_556_), .B(_550__bF_buf8), .C(_557_), .Y(_257__35_) );
	INVX1 INVX1_327 ( .A(bloque_in_1_36_), .Y(_558_) );
	OAI21X1 OAI21X1_470 ( .A(_550__bF_buf7), .B(RAM_entrada_94_), .C(reset_L_bF_buf38), .Y(_559_) );
	AOI21X1 AOI21X1_323 ( .A(_558_), .B(_550__bF_buf6), .C(_559_), .Y(_257__36_) );
	INVX1 INVX1_328 ( .A(bloque_in_1_37_), .Y(_560_) );
	OAI21X1 OAI21X1_471 ( .A(_550__bF_buf5), .B(RAM_entrada_93_), .C(reset_L_bF_buf37), .Y(_561_) );
	AOI21X1 AOI21X1_324 ( .A(_560_), .B(_550__bF_buf4), .C(_561_), .Y(_257__37_) );
	INVX1 INVX1_329 ( .A(bloque_in_1_38_), .Y(_562_) );
	OAI21X1 OAI21X1_472 ( .A(_550__bF_buf3), .B(RAM_entrada_95_), .C(reset_L_bF_buf36), .Y(_563_) );
	AOI21X1 AOI21X1_325 ( .A(_562_), .B(_550__bF_buf2), .C(_563_), .Y(_257__38_) );
	INVX1 INVX1_330 ( .A(bloque_in_1_39_), .Y(_564_) );
	OAI21X1 OAI21X1_473 ( .A(_550__bF_buf1), .B(RAM_entrada_95_), .C(reset_L_bF_buf35), .Y(_565_) );
	AOI21X1 AOI21X1_326 ( .A(_564_), .B(_550__bF_buf0), .C(_565_), .Y(_257__39_) );
	INVX1 INVX1_331 ( .A(bloque_in_1_40_), .Y(_566_) );
	OAI21X1 OAI21X1_474 ( .A(_550__bF_buf15), .B(RAM_entrada_86_), .C(reset_L_bF_buf34), .Y(_567_) );
	AOI21X1 AOI21X1_327 ( .A(_566_), .B(_550__bF_buf14), .C(_567_), .Y(_257__40_) );
	INVX1 INVX1_332 ( .A(bloque_in_1_41_), .Y(_568_) );
	OAI21X1 OAI21X1_475 ( .A(_550__bF_buf13), .B(RAM_entrada_84_bF_buf2), .C(reset_L_bF_buf33), .Y(_569_) );
	AOI21X1 AOI21X1_328 ( .A(_568_), .B(_550__bF_buf12), .C(_569_), .Y(_257__41_) );
	INVX1 INVX1_333 ( .A(bloque_in_1_42_), .Y(_570_) );
	OAI21X1 OAI21X1_476 ( .A(_550__bF_buf11), .B(RAM_entrada_77_), .C(reset_L_bF_buf32), .Y(_571_) );
	AOI21X1 AOI21X1_329 ( .A(_570_), .B(_550__bF_buf10), .C(_571_), .Y(_257__42_) );
	INVX1 INVX1_334 ( .A(bloque_in_1_43_), .Y(_572_) );
	OAI21X1 OAI21X1_477 ( .A(_550__bF_buf9), .B(RAM_entrada_46_), .C(reset_L_bF_buf31), .Y(_573_) );
	AOI21X1 AOI21X1_330 ( .A(_572_), .B(_550__bF_buf8), .C(_573_), .Y(_257__43_) );
	INVX1 INVX1_335 ( .A(bloque_in_1_44_), .Y(_574_) );
	OAI21X1 OAI21X1_478 ( .A(_550__bF_buf7), .B(RAM_entrada_82_), .C(reset_L_bF_buf30), .Y(_575_) );
	AOI21X1 AOI21X1_331 ( .A(_574_), .B(_550__bF_buf6), .C(_575_), .Y(_257__44_) );
	INVX1 INVX1_336 ( .A(bloque_in_1_45_), .Y(_576_) );
	OAI21X1 OAI21X1_479 ( .A(_550__bF_buf5), .B(RAM_entrada_92_), .C(reset_L_bF_buf29), .Y(_577_) );
	AOI21X1 AOI21X1_332 ( .A(_576_), .B(_550__bF_buf4), .C(_577_), .Y(_257__45_) );
	INVX1 INVX1_337 ( .A(bloque_in_1_46_), .Y(_578_) );
	OAI21X1 OAI21X1_480 ( .A(_550__bF_buf3), .B(RAM_entrada_71_bF_buf3), .C(reset_L_bF_buf28), .Y(_579_) );
	AOI21X1 AOI21X1_333 ( .A(_578_), .B(_550__bF_buf2), .C(_579_), .Y(_257__46_) );
	INVX1 INVX1_338 ( .A(bloque_in_1_47_), .Y(_580_) );
	OAI21X1 OAI21X1_481 ( .A(_550__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf27), .Y(_581_) );
	AOI21X1 AOI21X1_334 ( .A(_580_), .B(_550__bF_buf0), .C(_581_), .Y(_257__47_) );
	INVX1 INVX1_339 ( .A(bloque_in_1_48_), .Y(_582_) );
	OAI21X1 OAI21X1_482 ( .A(_550__bF_buf15), .B(RAM_entrada_92_), .C(reset_L_bF_buf26), .Y(_583_) );
	AOI21X1 AOI21X1_335 ( .A(_582_), .B(_550__bF_buf14), .C(_583_), .Y(_257__48_) );
	INVX1 INVX1_340 ( .A(bloque_in_1_49_), .Y(_584_) );
	OAI21X1 OAI21X1_483 ( .A(_550__bF_buf13), .B(RAM_entrada_84_bF_buf1), .C(reset_L_bF_buf25), .Y(_585_) );
	AOI21X1 AOI21X1_336 ( .A(_584_), .B(_550__bF_buf12), .C(_585_), .Y(_257__49_) );
	INVX1 INVX1_341 ( .A(bloque_in_1_50_), .Y(_586_) );
	OAI21X1 OAI21X1_484 ( .A(_550__bF_buf11), .B(RAM_entrada_86_), .C(reset_L_bF_buf24), .Y(_587_) );
	AOI21X1 AOI21X1_337 ( .A(_586_), .B(_550__bF_buf10), .C(_587_), .Y(_257__50_) );
	INVX1 INVX1_342 ( .A(bloque_in_1_51_), .Y(_588_) );
	OAI21X1 OAI21X1_485 ( .A(_550__bF_buf9), .B(RAM_entrada_86_), .C(reset_L_bF_buf23), .Y(_589_) );
	AOI21X1 AOI21X1_338 ( .A(_588_), .B(_550__bF_buf8), .C(_589_), .Y(_257__51_) );
	INVX1 INVX1_343 ( .A(bloque_in_1_52_), .Y(_590_) );
	OAI21X1 OAI21X1_486 ( .A(_550__bF_buf7), .B(vdd), .C(reset_L_bF_buf22), .Y(_591_) );
	AOI21X1 AOI21X1_339 ( .A(_590_), .B(_550__bF_buf6), .C(_591_), .Y(_257__52_) );
	INVX1 INVX1_344 ( .A(bloque_in_1_53_), .Y(_592_) );
	OAI21X1 OAI21X1_487 ( .A(_550__bF_buf5), .B(RAM_entrada_58_), .C(reset_L_bF_buf21), .Y(_593_) );
	AOI21X1 AOI21X1_340 ( .A(_592_), .B(_550__bF_buf4), .C(_593_), .Y(_257__53_) );
	INVX1 INVX1_345 ( .A(bloque_in_1_54_), .Y(_594_) );
	OAI21X1 OAI21X1_488 ( .A(_550__bF_buf3), .B(gnd), .C(reset_L_bF_buf20), .Y(_595_) );
	AOI21X1 AOI21X1_341 ( .A(_594_), .B(_550__bF_buf2), .C(_595_), .Y(_257__54_) );
	INVX1 INVX1_346 ( .A(bloque_in_1_55_), .Y(_596_) );
	OAI21X1 OAI21X1_489 ( .A(_550__bF_buf1), .B(RAM_entrada_71_bF_buf2), .C(reset_L_bF_buf19), .Y(_597_) );
	AOI21X1 AOI21X1_342 ( .A(_596_), .B(_550__bF_buf0), .C(_597_), .Y(_257__55_) );
	INVX1 INVX1_347 ( .A(bloque_in_1_56_), .Y(_598_) );
	OAI21X1 OAI21X1_490 ( .A(_550__bF_buf15), .B(RAM_entrada_88_), .C(reset_L_bF_buf18), .Y(_599_) );
	AOI21X1 AOI21X1_343 ( .A(_598_), .B(_550__bF_buf14), .C(_599_), .Y(_257__56_) );
	INVX1 INVX1_348 ( .A(bloque_in_1_57_), .Y(_600_) );
	OAI21X1 OAI21X1_491 ( .A(_550__bF_buf13), .B(RAM_entrada_93_), .C(reset_L_bF_buf17), .Y(_601_) );
	AOI21X1 AOI21X1_344 ( .A(_600_), .B(_550__bF_buf12), .C(_601_), .Y(_257__57_) );
	INVX1 INVX1_349 ( .A(bloque_in_1_58_), .Y(_602_) );
	OAI21X1 OAI21X1_492 ( .A(_550__bF_buf11), .B(RAM_entrada_58_), .C(reset_L_bF_buf16), .Y(_603_) );
	AOI21X1 AOI21X1_345 ( .A(_602_), .B(_550__bF_buf10), .C(_603_), .Y(_257__58_) );
	INVX1 INVX1_350 ( .A(bloque_in_1_59_), .Y(_604_) );
	OAI21X1 OAI21X1_493 ( .A(_550__bF_buf9), .B(RAM_entrada_85_), .C(reset_L_bF_buf15), .Y(_605_) );
	AOI21X1 AOI21X1_346 ( .A(_604_), .B(_550__bF_buf8), .C(_605_), .Y(_257__59_) );
	INVX1 INVX1_351 ( .A(bloque_in_1_60_), .Y(_606_) );
	OAI21X1 OAI21X1_494 ( .A(_550__bF_buf7), .B(RAM_entrada_71_bF_buf1), .C(reset_L_bF_buf14), .Y(_607_) );
	AOI21X1 AOI21X1_347 ( .A(_606_), .B(_550__bF_buf6), .C(_607_), .Y(_257__60_) );
	INVX1 INVX1_352 ( .A(bloque_in_1_61_), .Y(_608_) );
	OAI21X1 OAI21X1_495 ( .A(_550__bF_buf5), .B(RAM_entrada_93_), .C(reset_L_bF_buf13), .Y(_609_) );
	AOI21X1 AOI21X1_348 ( .A(_608_), .B(_550__bF_buf4), .C(_609_), .Y(_257__61_) );
	INVX1 INVX1_353 ( .A(bloque_in_1_62_), .Y(_610_) );
	OAI21X1 OAI21X1_496 ( .A(_550__bF_buf3), .B(RAM_entrada_84_bF_buf0), .C(reset_L_bF_buf12), .Y(_611_) );
	AOI21X1 AOI21X1_349 ( .A(_610_), .B(_550__bF_buf2), .C(_611_), .Y(_257__62_) );
	INVX1 INVX1_354 ( .A(bloque_in_1_63_), .Y(_612_) );
	OAI21X1 OAI21X1_497 ( .A(_550__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf11), .Y(_613_) );
	AOI21X1 AOI21X1_350 ( .A(_612_), .B(_550__bF_buf0), .C(_613_), .Y(_257__63_) );
	INVX1 INVX1_355 ( .A(bloque_in_1_64_), .Y(_614_) );
	OAI21X1 OAI21X1_498 ( .A(_550__bF_buf15), .B(RAM_entrada_71_bF_buf0), .C(reset_L_bF_buf10), .Y(_615_) );
	AOI21X1 AOI21X1_351 ( .A(_614_), .B(_550__bF_buf14), .C(_615_), .Y(_257__64_) );
	INVX1 INVX1_356 ( .A(bloque_in_1_65_), .Y(_616_) );
	OAI21X1 OAI21X1_499 ( .A(_550__bF_buf13), .B(RAM_entrada_95_), .C(reset_L_bF_buf9), .Y(_617_) );
	AOI21X1 AOI21X1_352 ( .A(_616_), .B(_550__bF_buf12), .C(_617_), .Y(_257__65_) );
	INVX1 INVX1_357 ( .A(bloque_in_1_66_), .Y(_618_) );
	OAI21X1 OAI21X1_500 ( .A(_550__bF_buf11), .B(RAM_entrada_92_), .C(reset_L_bF_buf8), .Y(_619_) );
	AOI21X1 AOI21X1_353 ( .A(_618_), .B(_550__bF_buf10), .C(_619_), .Y(_257__66_) );
	INVX1 INVX1_358 ( .A(bloque_in_1_67_), .Y(_620_) );
	OAI21X1 OAI21X1_501 ( .A(_550__bF_buf9), .B(RAM_entrada_92_), .C(reset_L_bF_buf7), .Y(_621_) );
	AOI21X1 AOI21X1_354 ( .A(_620_), .B(_550__bF_buf8), .C(_621_), .Y(_257__67_) );
	INVX1 INVX1_359 ( .A(bloque_in_1_68_), .Y(_622_) );
	OAI21X1 OAI21X1_502 ( .A(_550__bF_buf7), .B(RAM_entrada_71_bF_buf3), .C(reset_L_bF_buf6), .Y(_623_) );
	AOI21X1 AOI21X1_355 ( .A(_622_), .B(_550__bF_buf6), .C(_623_), .Y(_257__68_) );
	INVX1 INVX1_360 ( .A(bloque_in_1_69_), .Y(_624_) );
	OAI21X1 OAI21X1_503 ( .A(_550__bF_buf5), .B(RAM_entrada_84_bF_buf3), .C(reset_L_bF_buf5), .Y(_625_) );
	AOI21X1 AOI21X1_356 ( .A(_624_), .B(_550__bF_buf4), .C(_625_), .Y(_257__69_) );
	INVX1 INVX1_361 ( .A(bloque_in_1_70_), .Y(_626_) );
	OAI21X1 OAI21X1_504 ( .A(_550__bF_buf3), .B(RAM_entrada_84_bF_buf2), .C(reset_L_bF_buf4), .Y(_627_) );
	AOI21X1 AOI21X1_357 ( .A(_626_), .B(_550__bF_buf2), .C(_627_), .Y(_257__70_) );
	INVX1 INVX1_362 ( .A(bloque_in_1_71_), .Y(_628_) );
	OAI21X1 OAI21X1_505 ( .A(_550__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf3), .Y(_629_) );
	AOI21X1 AOI21X1_358 ( .A(_628_), .B(_550__bF_buf0), .C(_629_), .Y(_257__71_) );
	INVX1 INVX1_363 ( .A(bloque_in_1_72_), .Y(_630_) );
	OAI21X1 OAI21X1_506 ( .A(_550__bF_buf15), .B(RAM_entrada_89_), .C(reset_L_bF_buf2), .Y(_631_) );
	AOI21X1 AOI21X1_359 ( .A(_630_), .B(_550__bF_buf14), .C(_631_), .Y(_257__72_) );
	INVX1 INVX1_364 ( .A(bloque_in_1_73_), .Y(_632_) );
	OAI21X1 OAI21X1_507 ( .A(_550__bF_buf13), .B(RAM_entrada_82_), .C(reset_L_bF_buf1), .Y(_633_) );
	AOI21X1 AOI21X1_360 ( .A(_632_), .B(_550__bF_buf12), .C(_633_), .Y(_257__73_) );
	INVX1 INVX1_365 ( .A(bloque_in_1_74_), .Y(_634_) );
	OAI21X1 OAI21X1_508 ( .A(_550__bF_buf11), .B(RAM_entrada_92_), .C(reset_L_bF_buf0), .Y(_635_) );
	AOI21X1 AOI21X1_361 ( .A(_634_), .B(_550__bF_buf10), .C(_635_), .Y(_257__74_) );
	INVX1 INVX1_366 ( .A(bloque_in_1_75_), .Y(_636_) );
	OAI21X1 OAI21X1_509 ( .A(_550__bF_buf9), .B(RAM_entrada_85_), .C(reset_L_bF_buf49), .Y(_637_) );
	AOI21X1 AOI21X1_362 ( .A(_636_), .B(_550__bF_buf8), .C(_637_), .Y(_257__75_) );
	INVX1 INVX1_367 ( .A(bloque_in_1_76_), .Y(_638_) );
	OAI21X1 OAI21X1_510 ( .A(_550__bF_buf7), .B(RAM_entrada_82_), .C(reset_L_bF_buf48), .Y(_639_) );
	AOI21X1 AOI21X1_363 ( .A(_638_), .B(_550__bF_buf6), .C(_639_), .Y(_257__76_) );
	INVX1 INVX1_368 ( .A(bloque_in_1_77_), .Y(_640_) );
	OAI21X1 OAI21X1_511 ( .A(_550__bF_buf5), .B(RAM_entrada_46_), .C(reset_L_bF_buf47), .Y(_641_) );
	AOI21X1 AOI21X1_364 ( .A(_640_), .B(_550__bF_buf4), .C(_641_), .Y(_257__77_) );
	INVX1 INVX1_369 ( .A(bloque_in_1_78_), .Y(_642_) );
	OAI21X1 OAI21X1_512 ( .A(_550__bF_buf3), .B(RAM_entrada_46_), .C(reset_L_bF_buf46), .Y(_643_) );
	AOI21X1 AOI21X1_365 ( .A(_642_), .B(_550__bF_buf2), .C(_643_), .Y(_257__78_) );
	INVX1 INVX1_370 ( .A(bloque_in_1_79_), .Y(_644_) );
	OAI21X1 OAI21X1_513 ( .A(_550__bF_buf1), .B(vdd), .C(reset_L_bF_buf45), .Y(_645_) );
	AOI21X1 AOI21X1_366 ( .A(_644_), .B(_550__bF_buf0), .C(_645_), .Y(_257__79_) );
	INVX1 INVX1_371 ( .A(bloque_in_1_80_), .Y(_646_) );
	OAI21X1 OAI21X1_514 ( .A(_550__bF_buf15), .B(RAM_entrada_71_bF_buf2), .C(reset_L_bF_buf44), .Y(_647_) );
	AOI21X1 AOI21X1_367 ( .A(_646_), .B(_550__bF_buf14), .C(_647_), .Y(_257__80_) );
	INVX1 INVX1_372 ( .A(bloque_in_1_81_), .Y(_648_) );
	OAI21X1 OAI21X1_515 ( .A(_550__bF_buf13), .B(RAM_entrada_84_bF_buf1), .C(reset_L_bF_buf43), .Y(_649_) );
	AOI21X1 AOI21X1_368 ( .A(_648_), .B(_550__bF_buf12), .C(_649_), .Y(_257__81_) );
	INVX1 INVX1_373 ( .A(bloque_in_1_82_), .Y(_650_) );
	OAI21X1 OAI21X1_516 ( .A(_550__bF_buf11), .B(RAM_entrada_71_bF_buf1), .C(reset_L_bF_buf42), .Y(_651_) );
	AOI21X1 AOI21X1_369 ( .A(_650_), .B(_550__bF_buf10), .C(_651_), .Y(_257__82_) );
	INVX1 INVX1_374 ( .A(bloque_in_1_83_), .Y(_652_) );
	OAI21X1 OAI21X1_517 ( .A(_550__bF_buf9), .B(RAM_entrada_93_), .C(reset_L_bF_buf41), .Y(_653_) );
	AOI21X1 AOI21X1_370 ( .A(_652_), .B(_550__bF_buf8), .C(_653_), .Y(_257__83_) );
	INVX1 INVX1_375 ( .A(bloque_in_1_84_), .Y(_654_) );
	OAI21X1 OAI21X1_518 ( .A(_550__bF_buf7), .B(RAM_entrada_89_), .C(reset_L_bF_buf40), .Y(_655_) );
	AOI21X1 AOI21X1_371 ( .A(_654_), .B(_550__bF_buf6), .C(_655_), .Y(_257__84_) );
	INVX1 INVX1_376 ( .A(bloque_in_1_85_), .Y(_656_) );
	OAI21X1 OAI21X1_519 ( .A(_550__bF_buf5), .B(RAM_entrada_71_bF_buf0), .C(reset_L_bF_buf39), .Y(_657_) );
	AOI21X1 AOI21X1_372 ( .A(_656_), .B(_550__bF_buf4), .C(_657_), .Y(_257__85_) );
	INVX1 INVX1_377 ( .A(bloque_in_1_86_), .Y(_658_) );
	OAI21X1 OAI21X1_520 ( .A(_550__bF_buf3), .B(RAM_entrada_84_bF_buf0), .C(reset_L_bF_buf38), .Y(_659_) );
	AOI21X1 AOI21X1_373 ( .A(_658_), .B(_550__bF_buf2), .C(_659_), .Y(_257__86_) );
	INVX1 INVX1_378 ( .A(bloque_in_1_87_), .Y(_660_) );
	OAI21X1 OAI21X1_521 ( .A(_550__bF_buf1), .B(RAM_entrada_85_), .C(reset_L_bF_buf37), .Y(_661_) );
	AOI21X1 AOI21X1_374 ( .A(_660_), .B(_550__bF_buf0), .C(_661_), .Y(_257__87_) );
	INVX1 INVX1_379 ( .A(bloque_in_1_88_), .Y(_662_) );
	OAI21X1 OAI21X1_522 ( .A(_550__bF_buf15), .B(RAM_entrada_89_), .C(reset_L_bF_buf36), .Y(_663_) );
	AOI21X1 AOI21X1_375 ( .A(_662_), .B(_550__bF_buf14), .C(_663_), .Y(_257__88_) );
	INVX1 INVX1_380 ( .A(bloque_in_1_89_), .Y(_664_) );
	OAI21X1 OAI21X1_523 ( .A(_550__bF_buf13), .B(RAM_entrada_58_), .C(reset_L_bF_buf35), .Y(_665_) );
	AOI21X1 AOI21X1_376 ( .A(_664_), .B(_550__bF_buf12), .C(_665_), .Y(_257__89_) );
	INVX1 INVX1_381 ( .A(bloque_in_1_90_), .Y(_666_) );
	OAI21X1 OAI21X1_524 ( .A(_550__bF_buf11), .B(RAM_entrada_58_), .C(reset_L_bF_buf34), .Y(_667_) );
	AOI21X1 AOI21X1_377 ( .A(_666_), .B(_550__bF_buf10), .C(_667_), .Y(_257__90_) );
	INVX1 INVX1_382 ( .A(bloque_in_1_91_), .Y(_668_) );
	OAI21X1 OAI21X1_525 ( .A(_550__bF_buf9), .B(RAM_entrada_95_), .C(reset_L_bF_buf33), .Y(_669_) );
	AOI21X1 AOI21X1_378 ( .A(_668_), .B(_550__bF_buf8), .C(_669_), .Y(_257__91_) );
	INVX1 INVX1_383 ( .A(bloque_in_1_92_), .Y(_670_) );
	OAI21X1 OAI21X1_526 ( .A(_550__bF_buf7), .B(RAM_entrada_94_), .C(reset_L_bF_buf32), .Y(_671_) );
	AOI21X1 AOI21X1_379 ( .A(_670_), .B(_550__bF_buf6), .C(_671_), .Y(_257__92_) );
	INVX1 INVX1_384 ( .A(bloque_in_1_93_), .Y(_672_) );
	OAI21X1 OAI21X1_527 ( .A(_550__bF_buf5), .B(RAM_entrada_71_bF_buf3), .C(reset_L_bF_buf31), .Y(_673_) );
	AOI21X1 AOI21X1_380 ( .A(_672_), .B(_550__bF_buf4), .C(_673_), .Y(_257__93_) );
	INVX1 INVX1_385 ( .A(bloque_in_1_94_), .Y(_674_) );
	OAI21X1 OAI21X1_528 ( .A(_550__bF_buf3), .B(RAM_entrada_86_), .C(reset_L_bF_buf30), .Y(_675_) );
	AOI21X1 AOI21X1_381 ( .A(_674_), .B(_550__bF_buf2), .C(_675_), .Y(_257__94_) );
	INVX1 INVX1_386 ( .A(bloque_in_1_95_), .Y(_676_) );
	OAI21X1 OAI21X1_529 ( .A(_550__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf29), .Y(_677_) );
	AOI21X1 AOI21X1_382 ( .A(_676_), .B(_550__bF_buf0), .C(_677_), .Y(_257__95_) );
	INVX1 INVX1_387 ( .A(bloque_in_1_96_), .Y(_678_) );
	OAI21X1 OAI21X1_530 ( .A(_550__bF_buf15), .B(RAM_entrada_88_), .C(reset_L_bF_buf28), .Y(_679_) );
	AOI21X1 AOI21X1_383 ( .A(_678_), .B(_550__bF_buf14), .C(_679_), .Y(_257__96_) );
	INVX1 INVX1_388 ( .A(bloque_in_1_97_), .Y(_680_) );
	OAI21X1 OAI21X1_531 ( .A(_550__bF_buf13), .B(RAM_entrada_93_), .C(reset_L_bF_buf27), .Y(_681_) );
	AOI21X1 AOI21X1_384 ( .A(_680_), .B(_550__bF_buf12), .C(_681_), .Y(_257__97_) );
	INVX1 INVX1_389 ( .A(bloque_in_1_98_), .Y(_682_) );
	OAI21X1 OAI21X1_532 ( .A(_550__bF_buf11), .B(RAM_entrada_93_), .C(reset_L_bF_buf26), .Y(_683_) );
	AOI21X1 AOI21X1_385 ( .A(_682_), .B(_550__bF_buf10), .C(_683_), .Y(_257__98_) );
	INVX1 INVX1_390 ( .A(bloque_in_1_99_), .Y(_684_) );
	OAI21X1 OAI21X1_533 ( .A(_550__bF_buf9), .B(vdd), .C(reset_L_bF_buf25), .Y(_685_) );
	AOI21X1 AOI21X1_386 ( .A(_684_), .B(_550__bF_buf8), .C(_685_), .Y(_257__99_) );
	INVX1 INVX1_391 ( .A(bloque_in_1_100_), .Y(_686_) );
	OAI21X1 OAI21X1_534 ( .A(_550__bF_buf7), .B(RAM_entrada_89_), .C(reset_L_bF_buf24), .Y(_687_) );
	AOI21X1 AOI21X1_387 ( .A(_686_), .B(_550__bF_buf6), .C(_687_), .Y(_257__100_) );
	INVX1 INVX1_392 ( .A(bloque_in_1_101_), .Y(_688_) );
	OAI21X1 OAI21X1_535 ( .A(_550__bF_buf5), .B(RAM_entrada_82_), .C(reset_L_bF_buf23), .Y(_689_) );
	AOI21X1 AOI21X1_388 ( .A(_688_), .B(_550__bF_buf4), .C(_689_), .Y(_257__101_) );
	INVX1 INVX1_393 ( .A(bloque_in_1_102_), .Y(_690_) );
	OAI21X1 OAI21X1_536 ( .A(_550__bF_buf3), .B(RAM_entrada_71_bF_buf2), .C(reset_L_bF_buf22), .Y(_691_) );
	AOI21X1 AOI21X1_389 ( .A(_690_), .B(_550__bF_buf2), .C(_691_), .Y(_257__102_) );
	INVX1 INVX1_394 ( .A(bloque_in_1_103_), .Y(_692_) );
	OAI21X1 OAI21X1_537 ( .A(_550__bF_buf1), .B(RAM_entrada_71_bF_buf1), .C(reset_L_bF_buf21), .Y(_693_) );
	AOI21X1 AOI21X1_390 ( .A(_692_), .B(_550__bF_buf0), .C(_693_), .Y(_257__103_) );
	INVX1 INVX1_395 ( .A(bloque_in_1_104_), .Y(_694_) );
	OAI21X1 OAI21X1_538 ( .A(_550__bF_buf15), .B(RAM_entrada_92_), .C(reset_L_bF_buf20), .Y(_695_) );
	AOI21X1 AOI21X1_391 ( .A(_694_), .B(_550__bF_buf14), .C(_695_), .Y(_257__104_) );
	INVX1 INVX1_396 ( .A(bloque_in_1_105_), .Y(_696_) );
	OAI21X1 OAI21X1_539 ( .A(_550__bF_buf13), .B(RAM_entrada_88_), .C(reset_L_bF_buf19), .Y(_697_) );
	AOI21X1 AOI21X1_392 ( .A(_696_), .B(_550__bF_buf12), .C(_697_), .Y(_257__105_) );
	INVX1 INVX1_397 ( .A(bloque_in_1_106_), .Y(_698_) );
	OAI21X1 OAI21X1_540 ( .A(_550__bF_buf11), .B(RAM_entrada_88_), .C(reset_L_bF_buf18), .Y(_699_) );
	AOI21X1 AOI21X1_393 ( .A(_698_), .B(_550__bF_buf10), .C(_699_), .Y(_257__106_) );
	INVX1 INVX1_398 ( .A(bloque_in_1_107_), .Y(_700_) );
	OAI21X1 OAI21X1_541 ( .A(_550__bF_buf9), .B(vdd), .C(reset_L_bF_buf17), .Y(_701_) );
	AOI21X1 AOI21X1_394 ( .A(_700_), .B(_550__bF_buf8), .C(_701_), .Y(_257__107_) );
	INVX1 INVX1_399 ( .A(bloque_in_1_108_), .Y(_702_) );
	OAI21X1 OAI21X1_542 ( .A(_550__bF_buf7), .B(RAM_entrada_84_bF_buf3), .C(reset_L_bF_buf16), .Y(_703_) );
	AOI21X1 AOI21X1_395 ( .A(_702_), .B(_550__bF_buf6), .C(_703_), .Y(_257__108_) );
	INVX1 INVX1_400 ( .A(bloque_in_1_109_), .Y(_704_) );
	OAI21X1 OAI21X1_543 ( .A(_550__bF_buf5), .B(RAM_entrada_77_), .C(reset_L_bF_buf15), .Y(_705_) );
	AOI21X1 AOI21X1_396 ( .A(_704_), .B(_550__bF_buf4), .C(_705_), .Y(_257__109_) );
	INVX1 INVX1_401 ( .A(bloque_in_1_110_), .Y(_706_) );
	OAI21X1 OAI21X1_544 ( .A(_550__bF_buf3), .B(RAM_entrada_89_), .C(reset_L_bF_buf14), .Y(_707_) );
	AOI21X1 AOI21X1_397 ( .A(_706_), .B(_550__bF_buf2), .C(_707_), .Y(_257__110_) );
	INVX1 INVX1_402 ( .A(bloque_in_1_111_), .Y(_708_) );
	OAI21X1 OAI21X1_545 ( .A(_550__bF_buf1), .B(RAM_entrada_88_), .C(reset_L_bF_buf13), .Y(_709_) );
	AOI21X1 AOI21X1_398 ( .A(_708_), .B(_550__bF_buf0), .C(_709_), .Y(_257__111_) );
	INVX1 INVX1_403 ( .A(bloque_in_1_112_), .Y(_710_) );
	OAI21X1 OAI21X1_546 ( .A(_550__bF_buf15), .B(RAM_entrada_85_), .C(reset_L_bF_buf12), .Y(_711_) );
	AOI21X1 AOI21X1_399 ( .A(_710_), .B(_550__bF_buf14), .C(_711_), .Y(_257__112_) );
	INVX1 INVX1_404 ( .A(bloque_in_1_113_), .Y(_712_) );
	OAI21X1 OAI21X1_547 ( .A(_550__bF_buf13), .B(RAM_entrada_89_), .C(reset_L_bF_buf11), .Y(_713_) );
	AOI21X1 AOI21X1_400 ( .A(_712_), .B(_550__bF_buf12), .C(_713_), .Y(_257__113_) );
	INVX1 INVX1_405 ( .A(bloque_in_1_114_), .Y(_714_) );
	OAI21X1 OAI21X1_548 ( .A(_550__bF_buf11), .B(RAM_entrada_82_), .C(reset_L_bF_buf10), .Y(_715_) );
	AOI21X1 AOI21X1_401 ( .A(_714_), .B(_550__bF_buf10), .C(_715_), .Y(_257__114_) );
	INVX1 INVX1_406 ( .A(bloque_in_1_115_), .Y(_716_) );
	OAI21X1 OAI21X1_549 ( .A(_550__bF_buf9), .B(RAM_entrada_84_bF_buf2), .C(reset_L_bF_buf9), .Y(_717_) );
	AOI21X1 AOI21X1_402 ( .A(_716_), .B(_550__bF_buf8), .C(_717_), .Y(_257__115_) );
	INVX1 INVX1_407 ( .A(bloque_in_1_116_), .Y(_718_) );
	OAI21X1 OAI21X1_550 ( .A(_550__bF_buf7), .B(RAM_entrada_84_bF_buf1), .C(reset_L_bF_buf8), .Y(_719_) );
	AOI21X1 AOI21X1_403 ( .A(_718_), .B(_550__bF_buf6), .C(_719_), .Y(_257__116_) );
	INVX1 INVX1_408 ( .A(bloque_in_1_117_), .Y(_720_) );
	OAI21X1 OAI21X1_551 ( .A(_550__bF_buf5), .B(RAM_entrada_85_), .C(reset_L_bF_buf7), .Y(_721_) );
	AOI21X1 AOI21X1_404 ( .A(_720_), .B(_550__bF_buf4), .C(_721_), .Y(_257__117_) );
	INVX1 INVX1_409 ( .A(bloque_in_1_118_), .Y(_722_) );
	OAI21X1 OAI21X1_552 ( .A(_550__bF_buf3), .B(RAM_entrada_86_), .C(reset_L_bF_buf6), .Y(_723_) );
	AOI21X1 AOI21X1_405 ( .A(_722_), .B(_550__bF_buf2), .C(_723_), .Y(_257__118_) );
	INVX1 INVX1_410 ( .A(bloque_in_1_119_), .Y(_724_) );
	OAI21X1 OAI21X1_553 ( .A(_550__bF_buf1), .B(gnd), .C(reset_L_bF_buf5), .Y(_725_) );
	AOI21X1 AOI21X1_406 ( .A(_724_), .B(_550__bF_buf0), .C(_725_), .Y(_257__119_) );
	INVX1 INVX1_411 ( .A(bloque_in_1_120_), .Y(_726_) );
	OAI21X1 OAI21X1_554 ( .A(_550__bF_buf15), .B(RAM_entrada_88_), .C(reset_L_bF_buf4), .Y(_727_) );
	AOI21X1 AOI21X1_407 ( .A(_726_), .B(_550__bF_buf14), .C(_727_), .Y(_257__120_) );
	INVX1 INVX1_412 ( .A(bloque_in_1_121_), .Y(_728_) );
	OAI21X1 OAI21X1_555 ( .A(_550__bF_buf13), .B(RAM_entrada_89_), .C(reset_L_bF_buf3), .Y(_729_) );
	AOI21X1 AOI21X1_408 ( .A(_728_), .B(_550__bF_buf12), .C(_729_), .Y(_257__121_) );
	INVX1 INVX1_413 ( .A(bloque_in_1_122_), .Y(_730_) );
	OAI21X1 OAI21X1_556 ( .A(_550__bF_buf11), .B(RAM_entrada_94_), .C(reset_L_bF_buf2), .Y(_731_) );
	AOI21X1 AOI21X1_409 ( .A(_730_), .B(_550__bF_buf10), .C(_731_), .Y(_257__122_) );
	INVX1 INVX1_414 ( .A(bloque_in_1_123_), .Y(_732_) );
	OAI21X1 OAI21X1_557 ( .A(_550__bF_buf9), .B(vdd), .C(reset_L_bF_buf1), .Y(_733_) );
	AOI21X1 AOI21X1_410 ( .A(_732_), .B(_550__bF_buf8), .C(_733_), .Y(_257__123_) );
	INVX1 INVX1_415 ( .A(bloque_in_1_124_), .Y(_734_) );
	OAI21X1 OAI21X1_558 ( .A(_550__bF_buf7), .B(RAM_entrada_92_), .C(reset_L_bF_buf0), .Y(_735_) );
	AOI21X1 AOI21X1_411 ( .A(_734_), .B(_550__bF_buf6), .C(_735_), .Y(_257__124_) );
	INVX1 INVX1_416 ( .A(bloque_in_1_125_), .Y(_736_) );
	OAI21X1 OAI21X1_559 ( .A(_550__bF_buf5), .B(RAM_entrada_93_), .C(reset_L_bF_buf49), .Y(_737_) );
	AOI21X1 AOI21X1_412 ( .A(_736_), .B(_550__bF_buf4), .C(_737_), .Y(_257__125_) );
	INVX1 INVX1_417 ( .A(bloque_in_1_126_), .Y(_738_) );
	OAI21X1 OAI21X1_560 ( .A(_550__bF_buf3), .B(RAM_entrada_94_), .C(reset_L_bF_buf48), .Y(_739_) );
	AOI21X1 AOI21X1_413 ( .A(_738_), .B(_550__bF_buf2), .C(_739_), .Y(_257__126_) );
	INVX1 INVX1_418 ( .A(bloque_in_1_127_), .Y(_740_) );
	OAI21X1 OAI21X1_561 ( .A(_550__bF_buf1), .B(RAM_entrada_95_), .C(reset_L_bF_buf47), .Y(_741_) );
	AOI21X1 AOI21X1_414 ( .A(_740_), .B(_550__bF_buf0), .C(_741_), .Y(_257__127_) );
	INVX1 INVX1_419 ( .A(bloque_in_1_0_), .Y(_742_) );
	OAI21X1 OAI21X1_562 ( .A(_550__bF_buf15), .B(_2__0_), .C(reset_L_bF_buf46), .Y(_743_) );
	AOI21X1 AOI21X1_415 ( .A(_742_), .B(_550__bF_buf14), .C(_743_), .Y(_257__0_) );
	INVX1 INVX1_420 ( .A(bloque_in_1_1_), .Y(_744_) );
	OAI21X1 OAI21X1_563 ( .A(_550__bF_buf13), .B(_2__1_), .C(reset_L_bF_buf45), .Y(_745_) );
	AOI21X1 AOI21X1_416 ( .A(_744_), .B(_550__bF_buf12), .C(_745_), .Y(_257__1_) );
	INVX1 INVX1_421 ( .A(bloque_in_1_2_), .Y(_746_) );
	OAI21X1 OAI21X1_564 ( .A(_550__bF_buf11), .B(_2__2_), .C(reset_L_bF_buf44), .Y(_747_) );
	AOI21X1 AOI21X1_417 ( .A(_746_), .B(_550__bF_buf10), .C(_747_), .Y(_257__2_) );
	INVX1 INVX1_422 ( .A(bloque_in_1_3_), .Y(_748_) );
	OAI21X1 OAI21X1_565 ( .A(_550__bF_buf9), .B(_2__3_), .C(reset_L_bF_buf43), .Y(_749_) );
	AOI21X1 AOI21X1_418 ( .A(_748_), .B(_550__bF_buf8), .C(_749_), .Y(_257__3_) );
	INVX1 INVX1_423 ( .A(bloque_in_1_4_), .Y(_750_) );
	OAI21X1 OAI21X1_566 ( .A(_550__bF_buf7), .B(_2__4_), .C(reset_L_bF_buf42), .Y(_751_) );
	AOI21X1 AOI21X1_419 ( .A(_750_), .B(_550__bF_buf6), .C(_751_), .Y(_257__4_) );
	INVX1 INVX1_424 ( .A(bloque_in_1_5_), .Y(_752_) );
	OAI21X1 OAI21X1_567 ( .A(_550__bF_buf5), .B(_2__5_), .C(reset_L_bF_buf41), .Y(_753_) );
	AOI21X1 AOI21X1_420 ( .A(_752_), .B(_550__bF_buf4), .C(_753_), .Y(_257__5_) );
	INVX1 INVX1_425 ( .A(bloque_in_1_6_), .Y(_754_) );
	OAI21X1 OAI21X1_568 ( .A(_550__bF_buf3), .B(_2__6_), .C(reset_L_bF_buf40), .Y(_755_) );
	AOI21X1 AOI21X1_421 ( .A(_754_), .B(_550__bF_buf2), .C(_755_), .Y(_257__6_) );
	INVX1 INVX1_426 ( .A(bloque_in_1_7_), .Y(_756_) );
	OAI21X1 OAI21X1_569 ( .A(_550__bF_buf1), .B(_2__7_), .C(reset_L_bF_buf39), .Y(_757_) );
	AOI21X1 AOI21X1_422 ( .A(_756_), .B(_550__bF_buf0), .C(_757_), .Y(_257__7_) );
	INVX1 INVX1_427 ( .A(bloque_in_1_8_), .Y(_758_) );
	OAI21X1 OAI21X1_570 ( .A(_550__bF_buf15), .B(_2__8_), .C(reset_L_bF_buf38), .Y(_759_) );
	AOI21X1 AOI21X1_423 ( .A(_758_), .B(_550__bF_buf14), .C(_759_), .Y(_257__8_) );
	INVX1 INVX1_428 ( .A(bloque_in_1_9_), .Y(_760_) );
	OAI21X1 OAI21X1_571 ( .A(_550__bF_buf13), .B(_2__9_), .C(reset_L_bF_buf37), .Y(_761_) );
	AOI21X1 AOI21X1_424 ( .A(_760_), .B(_550__bF_buf12), .C(_761_), .Y(_257__9_) );
	INVX1 INVX1_429 ( .A(bloque_in_1_10_), .Y(_762_) );
	OAI21X1 OAI21X1_572 ( .A(_550__bF_buf11), .B(_2__10_), .C(reset_L_bF_buf36), .Y(_763_) );
	AOI21X1 AOI21X1_425 ( .A(_762_), .B(_550__bF_buf10), .C(_763_), .Y(_257__10_) );
	INVX1 INVX1_430 ( .A(bloque_in_1_11_), .Y(_764_) );
	OAI21X1 OAI21X1_573 ( .A(_550__bF_buf9), .B(_2__11_), .C(reset_L_bF_buf35), .Y(_765_) );
	AOI21X1 AOI21X1_426 ( .A(_764_), .B(_550__bF_buf8), .C(_765_), .Y(_257__11_) );
	INVX1 INVX1_431 ( .A(bloque_in_1_12_), .Y(_766_) );
	OAI21X1 OAI21X1_574 ( .A(_550__bF_buf7), .B(_2__12_), .C(reset_L_bF_buf34), .Y(_767_) );
	AOI21X1 AOI21X1_427 ( .A(_766_), .B(_550__bF_buf6), .C(_767_), .Y(_257__12_) );
	INVX1 INVX1_432 ( .A(bloque_in_1_13_), .Y(_768_) );
	OAI21X1 OAI21X1_575 ( .A(_550__bF_buf5), .B(_2__13_), .C(reset_L_bF_buf33), .Y(_769_) );
	AOI21X1 AOI21X1_428 ( .A(_768_), .B(_550__bF_buf4), .C(_769_), .Y(_257__13_) );
	INVX1 INVX1_433 ( .A(bloque_in_1_14_), .Y(_770_) );
	OAI21X1 OAI21X1_576 ( .A(_550__bF_buf3), .B(_2__14_), .C(reset_L_bF_buf32), .Y(_771_) );
	AOI21X1 AOI21X1_429 ( .A(_770_), .B(_550__bF_buf2), .C(_771_), .Y(_257__14_) );
	INVX1 INVX1_434 ( .A(bloque_in_1_15_), .Y(_772_) );
	OAI21X1 OAI21X1_577 ( .A(_550__bF_buf1), .B(_2__15_), .C(reset_L_bF_buf31), .Y(_773_) );
	AOI21X1 AOI21X1_430 ( .A(_772_), .B(_550__bF_buf0), .C(_773_), .Y(_257__15_) );
	INVX1 INVX1_435 ( .A(bloque_in_1_16_), .Y(_774_) );
	OAI21X1 OAI21X1_578 ( .A(_550__bF_buf15), .B(_2__16_), .C(reset_L_bF_buf30), .Y(_775_) );
	AOI21X1 AOI21X1_431 ( .A(_774_), .B(_550__bF_buf14), .C(_775_), .Y(_257__16_) );
	INVX1 INVX1_436 ( .A(bloque_in_1_17_), .Y(_776_) );
	OAI21X1 OAI21X1_579 ( .A(_550__bF_buf13), .B(_2__17_), .C(reset_L_bF_buf29), .Y(_777_) );
	AOI21X1 AOI21X1_432 ( .A(_776_), .B(_550__bF_buf12), .C(_777_), .Y(_257__17_) );
	INVX1 INVX1_437 ( .A(bloque_in_1_18_), .Y(_258_) );
	OAI21X1 OAI21X1_580 ( .A(_550__bF_buf11), .B(_2__18_), .C(reset_L_bF_buf28), .Y(_259_) );
	AOI21X1 AOI21X1_433 ( .A(_258_), .B(_550__bF_buf10), .C(_259_), .Y(_257__18_) );
	INVX1 INVX1_438 ( .A(bloque_in_1_19_), .Y(_260_) );
	OAI21X1 OAI21X1_581 ( .A(_550__bF_buf9), .B(_2__19_), .C(reset_L_bF_buf27), .Y(_261_) );
	AOI21X1 AOI21X1_434 ( .A(_260_), .B(_550__bF_buf8), .C(_261_), .Y(_257__19_) );
	INVX1 INVX1_439 ( .A(bloque_in_1_20_), .Y(_262_) );
	OAI21X1 OAI21X1_582 ( .A(_550__bF_buf7), .B(_2__20_), .C(reset_L_bF_buf26), .Y(_263_) );
	AOI21X1 AOI21X1_435 ( .A(_262_), .B(_550__bF_buf6), .C(_263_), .Y(_257__20_) );
	INVX1 INVX1_440 ( .A(bloque_in_1_21_), .Y(_264_) );
	OAI21X1 OAI21X1_583 ( .A(_550__bF_buf5), .B(_2__21_), .C(reset_L_bF_buf25), .Y(_265_) );
	AOI21X1 AOI21X1_436 ( .A(_264_), .B(_550__bF_buf4), .C(_265_), .Y(_257__21_) );
	INVX1 INVX1_441 ( .A(bloque_in_1_22_), .Y(_266_) );
	OAI21X1 OAI21X1_584 ( .A(_550__bF_buf3), .B(_2__22_), .C(reset_L_bF_buf24), .Y(_267_) );
	AOI21X1 AOI21X1_437 ( .A(_266_), .B(_550__bF_buf2), .C(_267_), .Y(_257__22_) );
	INVX1 INVX1_442 ( .A(bloque_in_1_23_), .Y(_268_) );
	OAI21X1 OAI21X1_585 ( .A(_550__bF_buf1), .B(_2__23_), .C(reset_L_bF_buf23), .Y(_269_) );
	AOI21X1 AOI21X1_438 ( .A(_268_), .B(_550__bF_buf0), .C(_269_), .Y(_257__23_) );
	INVX1 INVX1_443 ( .A(bloque_in_1_24_), .Y(_270_) );
	OAI21X1 OAI21X1_586 ( .A(_550__bF_buf15), .B(_2__24_), .C(reset_L_bF_buf22), .Y(_271_) );
	AOI21X1 AOI21X1_439 ( .A(_270_), .B(_550__bF_buf14), .C(_271_), .Y(_257__24_) );
	INVX1 INVX1_444 ( .A(bloque_in_1_25_), .Y(_272_) );
	OAI21X1 OAI21X1_587 ( .A(_550__bF_buf13), .B(_2__25_), .C(reset_L_bF_buf21), .Y(_273_) );
	AOI21X1 AOI21X1_440 ( .A(_272_), .B(_550__bF_buf12), .C(_273_), .Y(_257__25_) );
	INVX1 INVX1_445 ( .A(bloque_in_1_26_), .Y(_274_) );
	OAI21X1 OAI21X1_588 ( .A(_550__bF_buf11), .B(_2__26_), .C(reset_L_bF_buf20), .Y(_275_) );
	AOI21X1 AOI21X1_441 ( .A(_274_), .B(_550__bF_buf10), .C(_275_), .Y(_257__26_) );
	INVX1 INVX1_446 ( .A(bloque_in_1_27_), .Y(_276_) );
	OAI21X1 OAI21X1_589 ( .A(_550__bF_buf9), .B(_2__27_), .C(reset_L_bF_buf19), .Y(_277_) );
	AOI21X1 AOI21X1_442 ( .A(_276_), .B(_550__bF_buf8), .C(_277_), .Y(_257__27_) );
	INVX1 INVX1_447 ( .A(bloque_in_1_28_), .Y(_278_) );
	OAI21X1 OAI21X1_590 ( .A(_550__bF_buf7), .B(_2__28_), .C(reset_L_bF_buf18), .Y(_279_) );
	AOI21X1 AOI21X1_443 ( .A(_278_), .B(_550__bF_buf6), .C(_279_), .Y(_257__28_) );
	INVX1 INVX1_448 ( .A(bloque_in_1_29_), .Y(_280_) );
	OAI21X1 OAI21X1_591 ( .A(_550__bF_buf5), .B(_2__29_), .C(reset_L_bF_buf17), .Y(_281_) );
	AOI21X1 AOI21X1_444 ( .A(_280_), .B(_550__bF_buf4), .C(_281_), .Y(_257__29_) );
	INVX1 INVX1_449 ( .A(bloque_in_1_30_), .Y(_282_) );
	OAI21X1 OAI21X1_592 ( .A(_550__bF_buf3), .B(_2__30_), .C(reset_L_bF_buf16), .Y(_283_) );
	AOI21X1 AOI21X1_445 ( .A(_282_), .B(_550__bF_buf2), .C(_283_), .Y(_257__30_) );
	INVX1 INVX1_450 ( .A(bloque_in_1_31_), .Y(_284_) );
	OAI21X1 OAI21X1_593 ( .A(_550__bF_buf1), .B(_2__31_), .C(reset_L_bF_buf15), .Y(_285_) );
	AOI21X1 AOI21X1_446 ( .A(_284_), .B(_550__bF_buf0), .C(_285_), .Y(_257__31_) );
	INVX1 INVX1_451 ( .A(bloque_in_0_), .Y(_286_) );
	NOR2X1 NOR2X1_212 ( .A(concatenador_counter_1_bF_buf5), .B(concatenador_counter_0_bF_buf11), .Y(_287_) );
	NOR2X1 NOR2X1_213 ( .A(concatenador_counter_3_), .B(concatenador_counter_2_), .Y(_288_) );
	NOR2X1 NOR2X1_214 ( .A(concatenador_counter_5_), .B(concatenador_counter_4_), .Y(_289_) );
	NAND3X1 NAND3X1_122 ( .A(_287_), .B(_288_), .C(_289_), .Y(_290_) );
	OAI21X1 OAI21X1_594 ( .A(_290__bF_buf15), .B(_2__0_), .C(reset_L_bF_buf14), .Y(_291_) );
	AOI21X1 AOI21X1_447 ( .A(_286_), .B(_290__bF_buf14), .C(_291_), .Y(_256__0_) );
	INVX1 INVX1_452 ( .A(bloque_in_1_), .Y(_292_) );
	OAI21X1 OAI21X1_595 ( .A(_290__bF_buf13), .B(_2__1_), .C(reset_L_bF_buf13), .Y(_293_) );
	AOI21X1 AOI21X1_448 ( .A(_292_), .B(_290__bF_buf12), .C(_293_), .Y(_256__1_) );
	INVX1 INVX1_453 ( .A(bloque_in_2_), .Y(_294_) );
	OAI21X1 OAI21X1_596 ( .A(_290__bF_buf11), .B(_2__2_), .C(reset_L_bF_buf12), .Y(_295_) );
	AOI21X1 AOI21X1_449 ( .A(_294_), .B(_290__bF_buf10), .C(_295_), .Y(_256__2_) );
	INVX1 INVX1_454 ( .A(bloque_in_3_), .Y(_296_) );
	OAI21X1 OAI21X1_597 ( .A(_290__bF_buf9), .B(_2__3_), .C(reset_L_bF_buf11), .Y(_297_) );
	AOI21X1 AOI21X1_450 ( .A(_296_), .B(_290__bF_buf8), .C(_297_), .Y(_256__3_) );
	INVX1 INVX1_455 ( .A(bloque_in_4_), .Y(_298_) );
	OAI21X1 OAI21X1_598 ( .A(_290__bF_buf7), .B(_2__4_), .C(reset_L_bF_buf10), .Y(_299_) );
	AOI21X1 AOI21X1_451 ( .A(_298_), .B(_290__bF_buf6), .C(_299_), .Y(_256__4_) );
	INVX1 INVX1_456 ( .A(bloque_in_5_), .Y(_300_) );
	OAI21X1 OAI21X1_599 ( .A(_290__bF_buf5), .B(_2__5_), .C(reset_L_bF_buf9), .Y(_301_) );
	AOI21X1 AOI21X1_452 ( .A(_300_), .B(_290__bF_buf4), .C(_301_), .Y(_256__5_) );
	INVX1 INVX1_457 ( .A(bloque_in_6_), .Y(_302_) );
	OAI21X1 OAI21X1_600 ( .A(_290__bF_buf3), .B(_2__6_), .C(reset_L_bF_buf8), .Y(_303_) );
	AOI21X1 AOI21X1_453 ( .A(_302_), .B(_290__bF_buf2), .C(_303_), .Y(_256__6_) );
	INVX1 INVX1_458 ( .A(bloque_in_7_), .Y(_304_) );
	OAI21X1 OAI21X1_601 ( .A(_290__bF_buf1), .B(_2__7_), .C(reset_L_bF_buf7), .Y(_305_) );
	AOI21X1 AOI21X1_454 ( .A(_304_), .B(_290__bF_buf0), .C(_305_), .Y(_256__7_) );
	INVX1 INVX1_459 ( .A(bloque_in_8_), .Y(_306_) );
	OAI21X1 OAI21X1_602 ( .A(_290__bF_buf15), .B(_2__8_), .C(reset_L_bF_buf6), .Y(_307_) );
	AOI21X1 AOI21X1_455 ( .A(_306_), .B(_290__bF_buf14), .C(_307_), .Y(_256__8_) );
	INVX1 INVX1_460 ( .A(bloque_in_9_), .Y(_308_) );
	OAI21X1 OAI21X1_603 ( .A(_290__bF_buf13), .B(_2__9_), .C(reset_L_bF_buf5), .Y(_309_) );
	AOI21X1 AOI21X1_456 ( .A(_308_), .B(_290__bF_buf12), .C(_309_), .Y(_256__9_) );
	INVX1 INVX1_461 ( .A(bloque_in_10_), .Y(_310_) );
	OAI21X1 OAI21X1_604 ( .A(_290__bF_buf11), .B(_2__10_), .C(reset_L_bF_buf4), .Y(_311_) );
	AOI21X1 AOI21X1_457 ( .A(_310_), .B(_290__bF_buf10), .C(_311_), .Y(_256__10_) );
	INVX1 INVX1_462 ( .A(bloque_in_11_), .Y(_312_) );
	OAI21X1 OAI21X1_605 ( .A(_290__bF_buf9), .B(_2__11_), .C(reset_L_bF_buf3), .Y(_313_) );
	AOI21X1 AOI21X1_458 ( .A(_312_), .B(_290__bF_buf8), .C(_313_), .Y(_256__11_) );
	INVX1 INVX1_463 ( .A(bloque_in_12_), .Y(_314_) );
	OAI21X1 OAI21X1_606 ( .A(_290__bF_buf7), .B(_2__12_), .C(reset_L_bF_buf2), .Y(_315_) );
	AOI21X1 AOI21X1_459 ( .A(_314_), .B(_290__bF_buf6), .C(_315_), .Y(_256__12_) );
	INVX1 INVX1_464 ( .A(bloque_in_13_), .Y(_316_) );
	OAI21X1 OAI21X1_607 ( .A(_290__bF_buf5), .B(_2__13_), .C(reset_L_bF_buf1), .Y(_317_) );
	AOI21X1 AOI21X1_460 ( .A(_316_), .B(_290__bF_buf4), .C(_317_), .Y(_256__13_) );
	INVX1 INVX1_465 ( .A(bloque_in_14_), .Y(_318_) );
	OAI21X1 OAI21X1_608 ( .A(_290__bF_buf3), .B(_2__14_), .C(reset_L_bF_buf0), .Y(_319_) );
	AOI21X1 AOI21X1_461 ( .A(_318_), .B(_290__bF_buf2), .C(_319_), .Y(_256__14_) );
	INVX1 INVX1_466 ( .A(bloque_in_15_), .Y(_320_) );
	OAI21X1 OAI21X1_609 ( .A(_290__bF_buf1), .B(_2__15_), .C(reset_L_bF_buf49), .Y(_321_) );
	AOI21X1 AOI21X1_462 ( .A(_320_), .B(_290__bF_buf0), .C(_321_), .Y(_256__15_) );
	INVX1 INVX1_467 ( .A(bloque_in_16_), .Y(_322_) );
	OAI21X1 OAI21X1_610 ( .A(_290__bF_buf15), .B(_2__16_), .C(reset_L_bF_buf48), .Y(_323_) );
	AOI21X1 AOI21X1_463 ( .A(_322_), .B(_290__bF_buf14), .C(_323_), .Y(_256__16_) );
	INVX1 INVX1_468 ( .A(bloque_in_17_), .Y(_324_) );
	OAI21X1 OAI21X1_611 ( .A(_290__bF_buf13), .B(_2__17_), .C(reset_L_bF_buf47), .Y(_325_) );
	AOI21X1 AOI21X1_464 ( .A(_324_), .B(_290__bF_buf12), .C(_325_), .Y(_256__17_) );
	INVX1 INVX1_469 ( .A(bloque_in_18_), .Y(_326_) );
	OAI21X1 OAI21X1_612 ( .A(_290__bF_buf11), .B(_2__18_), .C(reset_L_bF_buf46), .Y(_327_) );
	AOI21X1 AOI21X1_465 ( .A(_326_), .B(_290__bF_buf10), .C(_327_), .Y(_256__18_) );
	INVX1 INVX1_470 ( .A(bloque_in_19_), .Y(_328_) );
	OAI21X1 OAI21X1_613 ( .A(_290__bF_buf9), .B(_2__19_), .C(reset_L_bF_buf45), .Y(_329_) );
	AOI21X1 AOI21X1_466 ( .A(_328_), .B(_290__bF_buf8), .C(_329_), .Y(_256__19_) );
	INVX1 INVX1_471 ( .A(bloque_in_20_), .Y(_330_) );
	OAI21X1 OAI21X1_614 ( .A(_290__bF_buf7), .B(_2__20_), .C(reset_L_bF_buf44), .Y(_331_) );
	AOI21X1 AOI21X1_467 ( .A(_330_), .B(_290__bF_buf6), .C(_331_), .Y(_256__20_) );
	INVX1 INVX1_472 ( .A(bloque_in_21_), .Y(_332_) );
	OAI21X1 OAI21X1_615 ( .A(_290__bF_buf5), .B(_2__21_), .C(reset_L_bF_buf43), .Y(_333_) );
	AOI21X1 AOI21X1_468 ( .A(_332_), .B(_290__bF_buf4), .C(_333_), .Y(_256__21_) );
	INVX1 INVX1_473 ( .A(bloque_in_22_), .Y(_334_) );
	OAI21X1 OAI21X1_616 ( .A(_290__bF_buf3), .B(_2__22_), .C(reset_L_bF_buf42), .Y(_335_) );
	AOI21X1 AOI21X1_469 ( .A(_334_), .B(_290__bF_buf2), .C(_335_), .Y(_256__22_) );
	INVX1 INVX1_474 ( .A(bloque_in_23_), .Y(_336_) );
	OAI21X1 OAI21X1_617 ( .A(_290__bF_buf1), .B(_2__23_), .C(reset_L_bF_buf41), .Y(_337_) );
	AOI21X1 AOI21X1_470 ( .A(_336_), .B(_290__bF_buf0), .C(_337_), .Y(_256__23_) );
	INVX1 INVX1_475 ( .A(bloque_in_24_), .Y(_338_) );
	OAI21X1 OAI21X1_618 ( .A(_290__bF_buf15), .B(_2__24_), .C(reset_L_bF_buf40), .Y(_339_) );
	AOI21X1 AOI21X1_471 ( .A(_338_), .B(_290__bF_buf14), .C(_339_), .Y(_256__24_) );
	INVX1 INVX1_476 ( .A(bloque_in_25_), .Y(_340_) );
	OAI21X1 OAI21X1_619 ( .A(_290__bF_buf13), .B(_2__25_), .C(reset_L_bF_buf39), .Y(_341_) );
	AOI21X1 AOI21X1_472 ( .A(_340_), .B(_290__bF_buf12), .C(_341_), .Y(_256__25_) );
	INVX1 INVX1_477 ( .A(bloque_in_26_), .Y(_342_) );
	OAI21X1 OAI21X1_620 ( .A(_290__bF_buf11), .B(_2__26_), .C(reset_L_bF_buf38), .Y(_343_) );
	AOI21X1 AOI21X1_473 ( .A(_342_), .B(_290__bF_buf10), .C(_343_), .Y(_256__26_) );
	INVX1 INVX1_478 ( .A(bloque_in_27_), .Y(_344_) );
	OAI21X1 OAI21X1_621 ( .A(_290__bF_buf9), .B(_2__27_), .C(reset_L_bF_buf37), .Y(_345_) );
	AOI21X1 AOI21X1_474 ( .A(_344_), .B(_290__bF_buf8), .C(_345_), .Y(_256__27_) );
	INVX1 INVX1_479 ( .A(bloque_in_28_), .Y(_346_) );
	OAI21X1 OAI21X1_622 ( .A(_290__bF_buf7), .B(_2__28_), .C(reset_L_bF_buf36), .Y(_347_) );
	AOI21X1 AOI21X1_475 ( .A(_346_), .B(_290__bF_buf6), .C(_347_), .Y(_256__28_) );
	INVX1 INVX1_480 ( .A(bloque_in_29_), .Y(_348_) );
	OAI21X1 OAI21X1_623 ( .A(_290__bF_buf5), .B(_2__29_), .C(reset_L_bF_buf35), .Y(_349_) );
	AOI21X1 AOI21X1_476 ( .A(_348_), .B(_290__bF_buf4), .C(_349_), .Y(_256__29_) );
	INVX1 INVX1_481 ( .A(bloque_in_30_), .Y(_350_) );
	OAI21X1 OAI21X1_624 ( .A(_290__bF_buf3), .B(_2__30_), .C(reset_L_bF_buf34), .Y(_351_) );
	AOI21X1 AOI21X1_477 ( .A(_350_), .B(_290__bF_buf2), .C(_351_), .Y(_256__30_) );
	INVX1 INVX1_482 ( .A(bloque_in_31_), .Y(_352_) );
	OAI21X1 OAI21X1_625 ( .A(_290__bF_buf1), .B(_2__31_), .C(reset_L_bF_buf33), .Y(_353_) );
	AOI21X1 AOI21X1_478 ( .A(_352_), .B(_290__bF_buf0), .C(_353_), .Y(_256__31_) );
	INVX1 INVX1_483 ( .A(bloque_in_32_), .Y(_354_) );
	OAI21X1 OAI21X1_626 ( .A(_290__bF_buf15), .B(RAM_entrada_89_), .C(reset_L_bF_buf32), .Y(_355_) );
	AOI21X1 AOI21X1_479 ( .A(_354_), .B(_290__bF_buf14), .C(_355_), .Y(_256__32_) );
	INVX1 INVX1_484 ( .A(bloque_in_33_), .Y(_356_) );
	OAI21X1 OAI21X1_627 ( .A(_290__bF_buf13), .B(RAM_entrada_77_), .C(reset_L_bF_buf31), .Y(_357_) );
	AOI21X1 AOI21X1_480 ( .A(_356_), .B(_290__bF_buf12), .C(_357_), .Y(_256__33_) );
	INVX1 INVX1_485 ( .A(bloque_in_34_), .Y(_358_) );
	OAI21X1 OAI21X1_628 ( .A(_290__bF_buf11), .B(RAM_entrada_84_bF_buf0), .C(reset_L_bF_buf30), .Y(_359_) );
	AOI21X1 AOI21X1_481 ( .A(_358_), .B(_290__bF_buf10), .C(_359_), .Y(_256__34_) );
	INVX1 INVX1_486 ( .A(bloque_in_35_), .Y(_360_) );
	OAI21X1 OAI21X1_629 ( .A(_290__bF_buf9), .B(RAM_entrada_94_), .C(reset_L_bF_buf29), .Y(_361_) );
	AOI21X1 AOI21X1_482 ( .A(_360_), .B(_290__bF_buf8), .C(_361_), .Y(_256__35_) );
	INVX1 INVX1_487 ( .A(bloque_in_36_), .Y(_362_) );
	OAI21X1 OAI21X1_630 ( .A(_290__bF_buf7), .B(RAM_entrada_94_), .C(reset_L_bF_buf28), .Y(_363_) );
	AOI21X1 AOI21X1_483 ( .A(_362_), .B(_290__bF_buf6), .C(_363_), .Y(_256__36_) );
	INVX1 INVX1_488 ( .A(bloque_in_37_), .Y(_364_) );
	OAI21X1 OAI21X1_631 ( .A(_290__bF_buf5), .B(RAM_entrada_93_), .C(reset_L_bF_buf27), .Y(_365_) );
	AOI21X1 AOI21X1_484 ( .A(_364_), .B(_290__bF_buf4), .C(_365_), .Y(_256__37_) );
	INVX1 INVX1_489 ( .A(bloque_in_38_), .Y(_366_) );
	OAI21X1 OAI21X1_632 ( .A(_290__bF_buf3), .B(RAM_entrada_95_), .C(reset_L_bF_buf26), .Y(_367_) );
	AOI21X1 AOI21X1_485 ( .A(_366_), .B(_290__bF_buf2), .C(_367_), .Y(_256__38_) );
	INVX1 INVX1_490 ( .A(bloque_in_39_), .Y(_368_) );
	OAI21X1 OAI21X1_633 ( .A(_290__bF_buf1), .B(RAM_entrada_95_), .C(reset_L_bF_buf25), .Y(_369_) );
	AOI21X1 AOI21X1_486 ( .A(_368_), .B(_290__bF_buf0), .C(_369_), .Y(_256__39_) );
	INVX1 INVX1_491 ( .A(bloque_in_40_), .Y(_370_) );
	OAI21X1 OAI21X1_634 ( .A(_290__bF_buf15), .B(RAM_entrada_86_), .C(reset_L_bF_buf24), .Y(_371_) );
	AOI21X1 AOI21X1_487 ( .A(_370_), .B(_290__bF_buf14), .C(_371_), .Y(_256__40_) );
	INVX1 INVX1_492 ( .A(bloque_in_41_), .Y(_372_) );
	OAI21X1 OAI21X1_635 ( .A(_290__bF_buf13), .B(RAM_entrada_84_bF_buf3), .C(reset_L_bF_buf23), .Y(_373_) );
	AOI21X1 AOI21X1_488 ( .A(_372_), .B(_290__bF_buf12), .C(_373_), .Y(_256__41_) );
	INVX1 INVX1_493 ( .A(bloque_in_42_), .Y(_374_) );
	OAI21X1 OAI21X1_636 ( .A(_290__bF_buf11), .B(RAM_entrada_77_), .C(reset_L_bF_buf22), .Y(_375_) );
	AOI21X1 AOI21X1_489 ( .A(_374_), .B(_290__bF_buf10), .C(_375_), .Y(_256__42_) );
	INVX1 INVX1_494 ( .A(bloque_in_43_), .Y(_376_) );
	OAI21X1 OAI21X1_637 ( .A(_290__bF_buf9), .B(RAM_entrada_46_), .C(reset_L_bF_buf21), .Y(_377_) );
	AOI21X1 AOI21X1_490 ( .A(_376_), .B(_290__bF_buf8), .C(_377_), .Y(_256__43_) );
	INVX1 INVX1_495 ( .A(bloque_in_44_), .Y(_378_) );
	OAI21X1 OAI21X1_638 ( .A(_290__bF_buf7), .B(RAM_entrada_82_), .C(reset_L_bF_buf20), .Y(_379_) );
	AOI21X1 AOI21X1_491 ( .A(_378_), .B(_290__bF_buf6), .C(_379_), .Y(_256__44_) );
	INVX1 INVX1_496 ( .A(bloque_in_45_), .Y(_380_) );
	OAI21X1 OAI21X1_639 ( .A(_290__bF_buf5), .B(RAM_entrada_92_), .C(reset_L_bF_buf19), .Y(_381_) );
	AOI21X1 AOI21X1_492 ( .A(_380_), .B(_290__bF_buf4), .C(_381_), .Y(_256__45_) );
	INVX1 INVX1_497 ( .A(bloque_in_46_), .Y(_382_) );
	OAI21X1 OAI21X1_640 ( .A(_290__bF_buf3), .B(RAM_entrada_71_bF_buf0), .C(reset_L_bF_buf18), .Y(_383_) );
	AOI21X1 AOI21X1_493 ( .A(_382_), .B(_290__bF_buf2), .C(_383_), .Y(_256__46_) );
	INVX1 INVX1_498 ( .A(bloque_in_47_), .Y(_384_) );
	OAI21X1 OAI21X1_641 ( .A(_290__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf17), .Y(_385_) );
	AOI21X1 AOI21X1_494 ( .A(_384_), .B(_290__bF_buf0), .C(_385_), .Y(_256__47_) );
	INVX1 INVX1_499 ( .A(bloque_in_48_), .Y(_386_) );
	OAI21X1 OAI21X1_642 ( .A(_290__bF_buf15), .B(RAM_entrada_92_), .C(reset_L_bF_buf16), .Y(_387_) );
	AOI21X1 AOI21X1_495 ( .A(_386_), .B(_290__bF_buf14), .C(_387_), .Y(_256__48_) );
	INVX1 INVX1_500 ( .A(bloque_in_49_), .Y(_388_) );
	OAI21X1 OAI21X1_643 ( .A(_290__bF_buf13), .B(RAM_entrada_84_bF_buf2), .C(reset_L_bF_buf15), .Y(_389_) );
	AOI21X1 AOI21X1_496 ( .A(_388_), .B(_290__bF_buf12), .C(_389_), .Y(_256__49_) );
	INVX1 INVX1_501 ( .A(bloque_in_50_), .Y(_390_) );
	OAI21X1 OAI21X1_644 ( .A(_290__bF_buf11), .B(RAM_entrada_86_), .C(reset_L_bF_buf14), .Y(_391_) );
	AOI21X1 AOI21X1_497 ( .A(_390_), .B(_290__bF_buf10), .C(_391_), .Y(_256__50_) );
	INVX1 INVX1_502 ( .A(bloque_in_51_), .Y(_392_) );
	OAI21X1 OAI21X1_645 ( .A(_290__bF_buf9), .B(RAM_entrada_86_), .C(reset_L_bF_buf13), .Y(_393_) );
	AOI21X1 AOI21X1_498 ( .A(_392_), .B(_290__bF_buf8), .C(_393_), .Y(_256__51_) );
	INVX1 INVX1_503 ( .A(bloque_in_52_), .Y(_394_) );
	OAI21X1 OAI21X1_646 ( .A(_290__bF_buf7), .B(vdd), .C(reset_L_bF_buf12), .Y(_395_) );
	AOI21X1 AOI21X1_499 ( .A(_394_), .B(_290__bF_buf6), .C(_395_), .Y(_256__52_) );
	INVX1 INVX1_504 ( .A(bloque_in_53_), .Y(_396_) );
	OAI21X1 OAI21X1_647 ( .A(_290__bF_buf5), .B(RAM_entrada_58_), .C(reset_L_bF_buf11), .Y(_397_) );
	AOI21X1 AOI21X1_500 ( .A(_396_), .B(_290__bF_buf4), .C(_397_), .Y(_256__53_) );
	INVX1 INVX1_505 ( .A(bloque_in_54_), .Y(_398_) );
	OAI21X1 OAI21X1_648 ( .A(_290__bF_buf3), .B(gnd), .C(reset_L_bF_buf10), .Y(_399_) );
	AOI21X1 AOI21X1_501 ( .A(_398_), .B(_290__bF_buf2), .C(_399_), .Y(_256__54_) );
	INVX1 INVX1_506 ( .A(bloque_in_55_), .Y(_400_) );
	OAI21X1 OAI21X1_649 ( .A(_290__bF_buf1), .B(RAM_entrada_71_bF_buf3), .C(reset_L_bF_buf9), .Y(_401_) );
	AOI21X1 AOI21X1_502 ( .A(_400_), .B(_290__bF_buf0), .C(_401_), .Y(_256__55_) );
	INVX1 INVX1_507 ( .A(bloque_in_56_), .Y(_402_) );
	OAI21X1 OAI21X1_650 ( .A(_290__bF_buf15), .B(RAM_entrada_88_), .C(reset_L_bF_buf8), .Y(_403_) );
	AOI21X1 AOI21X1_503 ( .A(_402_), .B(_290__bF_buf14), .C(_403_), .Y(_256__56_) );
	INVX1 INVX1_508 ( .A(bloque_in_57_), .Y(_404_) );
	OAI21X1 OAI21X1_651 ( .A(_290__bF_buf13), .B(RAM_entrada_93_), .C(reset_L_bF_buf7), .Y(_405_) );
	AOI21X1 AOI21X1_504 ( .A(_404_), .B(_290__bF_buf12), .C(_405_), .Y(_256__57_) );
	INVX1 INVX1_509 ( .A(bloque_in_58_), .Y(_406_) );
	OAI21X1 OAI21X1_652 ( .A(_290__bF_buf11), .B(RAM_entrada_58_), .C(reset_L_bF_buf6), .Y(_407_) );
	AOI21X1 AOI21X1_505 ( .A(_406_), .B(_290__bF_buf10), .C(_407_), .Y(_256__58_) );
	INVX1 INVX1_510 ( .A(bloque_in_59_), .Y(_408_) );
	OAI21X1 OAI21X1_653 ( .A(_290__bF_buf9), .B(RAM_entrada_85_), .C(reset_L_bF_buf5), .Y(_409_) );
	AOI21X1 AOI21X1_506 ( .A(_408_), .B(_290__bF_buf8), .C(_409_), .Y(_256__59_) );
	INVX1 INVX1_511 ( .A(bloque_in_60_), .Y(_410_) );
	OAI21X1 OAI21X1_654 ( .A(_290__bF_buf7), .B(RAM_entrada_71_bF_buf2), .C(reset_L_bF_buf4), .Y(_411_) );
	AOI21X1 AOI21X1_507 ( .A(_410_), .B(_290__bF_buf6), .C(_411_), .Y(_256__60_) );
	INVX1 INVX1_512 ( .A(bloque_in_61_), .Y(_412_) );
	OAI21X1 OAI21X1_655 ( .A(_290__bF_buf5), .B(RAM_entrada_93_), .C(reset_L_bF_buf3), .Y(_413_) );
	AOI21X1 AOI21X1_508 ( .A(_412_), .B(_290__bF_buf4), .C(_413_), .Y(_256__61_) );
	INVX1 INVX1_513 ( .A(bloque_in_62_), .Y(_414_) );
	OAI21X1 OAI21X1_656 ( .A(_290__bF_buf3), .B(RAM_entrada_84_bF_buf1), .C(reset_L_bF_buf2), .Y(_415_) );
	AOI21X1 AOI21X1_509 ( .A(_414_), .B(_290__bF_buf2), .C(_415_), .Y(_256__62_) );
	INVX1 INVX1_514 ( .A(bloque_in_63_), .Y(_416_) );
	OAI21X1 OAI21X1_657 ( .A(_290__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf1), .Y(_417_) );
	AOI21X1 AOI21X1_510 ( .A(_416_), .B(_290__bF_buf0), .C(_417_), .Y(_256__63_) );
	INVX1 INVX1_515 ( .A(bloque_in_64_), .Y(_418_) );
	OAI21X1 OAI21X1_658 ( .A(_290__bF_buf15), .B(RAM_entrada_71_bF_buf1), .C(reset_L_bF_buf0), .Y(_419_) );
	AOI21X1 AOI21X1_511 ( .A(_418_), .B(_290__bF_buf14), .C(_419_), .Y(_256__64_) );
	INVX1 INVX1_516 ( .A(bloque_in_65_), .Y(_420_) );
	OAI21X1 OAI21X1_659 ( .A(_290__bF_buf13), .B(RAM_entrada_95_), .C(reset_L_bF_buf49), .Y(_421_) );
	AOI21X1 AOI21X1_512 ( .A(_420_), .B(_290__bF_buf12), .C(_421_), .Y(_256__65_) );
	INVX1 INVX1_517 ( .A(bloque_in_66_), .Y(_422_) );
	OAI21X1 OAI21X1_660 ( .A(_290__bF_buf11), .B(RAM_entrada_92_), .C(reset_L_bF_buf48), .Y(_423_) );
	AOI21X1 AOI21X1_513 ( .A(_422_), .B(_290__bF_buf10), .C(_423_), .Y(_256__66_) );
	INVX1 INVX1_518 ( .A(bloque_in_67_), .Y(_424_) );
	OAI21X1 OAI21X1_661 ( .A(_290__bF_buf9), .B(RAM_entrada_92_), .C(reset_L_bF_buf47), .Y(_425_) );
	AOI21X1 AOI21X1_514 ( .A(_424_), .B(_290__bF_buf8), .C(_425_), .Y(_256__67_) );
	INVX1 INVX1_519 ( .A(bloque_in_68_), .Y(_426_) );
	OAI21X1 OAI21X1_662 ( .A(_290__bF_buf7), .B(RAM_entrada_71_bF_buf0), .C(reset_L_bF_buf46), .Y(_427_) );
	AOI21X1 AOI21X1_515 ( .A(_426_), .B(_290__bF_buf6), .C(_427_), .Y(_256__68_) );
	INVX1 INVX1_520 ( .A(bloque_in_69_), .Y(_428_) );
	OAI21X1 OAI21X1_663 ( .A(_290__bF_buf5), .B(RAM_entrada_84_bF_buf0), .C(reset_L_bF_buf45), .Y(_429_) );
	AOI21X1 AOI21X1_516 ( .A(_428_), .B(_290__bF_buf4), .C(_429_), .Y(_256__69_) );
	INVX1 INVX1_521 ( .A(bloque_in_70_), .Y(_430_) );
	OAI21X1 OAI21X1_664 ( .A(_290__bF_buf3), .B(RAM_entrada_84_bF_buf3), .C(reset_L_bF_buf44), .Y(_431_) );
	AOI21X1 AOI21X1_517 ( .A(_430_), .B(_290__bF_buf2), .C(_431_), .Y(_256__70_) );
	INVX1 INVX1_522 ( .A(bloque_in_71_), .Y(_432_) );
	OAI21X1 OAI21X1_665 ( .A(_290__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf43), .Y(_433_) );
	AOI21X1 AOI21X1_518 ( .A(_432_), .B(_290__bF_buf0), .C(_433_), .Y(_256__71_) );
	INVX1 INVX1_523 ( .A(bloque_in_72_), .Y(_434_) );
	OAI21X1 OAI21X1_666 ( .A(_290__bF_buf15), .B(RAM_entrada_89_), .C(reset_L_bF_buf42), .Y(_435_) );
	AOI21X1 AOI21X1_519 ( .A(_434_), .B(_290__bF_buf14), .C(_435_), .Y(_256__72_) );
	INVX1 INVX1_524 ( .A(bloque_in_73_), .Y(_436_) );
	OAI21X1 OAI21X1_667 ( .A(_290__bF_buf13), .B(RAM_entrada_82_), .C(reset_L_bF_buf41), .Y(_437_) );
	AOI21X1 AOI21X1_520 ( .A(_436_), .B(_290__bF_buf12), .C(_437_), .Y(_256__73_) );
	INVX1 INVX1_525 ( .A(bloque_in_74_), .Y(_438_) );
	OAI21X1 OAI21X1_668 ( .A(_290__bF_buf11), .B(RAM_entrada_92_), .C(reset_L_bF_buf40), .Y(_439_) );
	AOI21X1 AOI21X1_521 ( .A(_438_), .B(_290__bF_buf10), .C(_439_), .Y(_256__74_) );
	INVX1 INVX1_526 ( .A(bloque_in_75_), .Y(_440_) );
	OAI21X1 OAI21X1_669 ( .A(_290__bF_buf9), .B(RAM_entrada_85_), .C(reset_L_bF_buf39), .Y(_441_) );
	AOI21X1 AOI21X1_522 ( .A(_440_), .B(_290__bF_buf8), .C(_441_), .Y(_256__75_) );
	INVX1 INVX1_527 ( .A(bloque_in_76_), .Y(_442_) );
	OAI21X1 OAI21X1_670 ( .A(_290__bF_buf7), .B(RAM_entrada_82_), .C(reset_L_bF_buf38), .Y(_443_) );
	AOI21X1 AOI21X1_523 ( .A(_442_), .B(_290__bF_buf6), .C(_443_), .Y(_256__76_) );
	INVX1 INVX1_528 ( .A(bloque_in_77_), .Y(_444_) );
	OAI21X1 OAI21X1_671 ( .A(_290__bF_buf5), .B(RAM_entrada_46_), .C(reset_L_bF_buf37), .Y(_445_) );
	AOI21X1 AOI21X1_524 ( .A(_444_), .B(_290__bF_buf4), .C(_445_), .Y(_256__77_) );
	INVX1 INVX1_529 ( .A(bloque_in_78_), .Y(_446_) );
	OAI21X1 OAI21X1_672 ( .A(_290__bF_buf3), .B(RAM_entrada_46_), .C(reset_L_bF_buf36), .Y(_447_) );
	AOI21X1 AOI21X1_525 ( .A(_446_), .B(_290__bF_buf2), .C(_447_), .Y(_256__78_) );
	INVX1 INVX1_530 ( .A(bloque_in_79_), .Y(_448_) );
	OAI21X1 OAI21X1_673 ( .A(_290__bF_buf1), .B(vdd), .C(reset_L_bF_buf35), .Y(_449_) );
	AOI21X1 AOI21X1_526 ( .A(_448_), .B(_290__bF_buf0), .C(_449_), .Y(_256__79_) );
	INVX1 INVX1_531 ( .A(bloque_in_80_), .Y(_450_) );
	OAI21X1 OAI21X1_674 ( .A(_290__bF_buf15), .B(RAM_entrada_71_bF_buf3), .C(reset_L_bF_buf34), .Y(_451_) );
	AOI21X1 AOI21X1_527 ( .A(_450_), .B(_290__bF_buf14), .C(_451_), .Y(_256__80_) );
	INVX1 INVX1_532 ( .A(bloque_in_81_), .Y(_452_) );
	OAI21X1 OAI21X1_675 ( .A(_290__bF_buf13), .B(RAM_entrada_84_bF_buf2), .C(reset_L_bF_buf33), .Y(_453_) );
	AOI21X1 AOI21X1_528 ( .A(_452_), .B(_290__bF_buf12), .C(_453_), .Y(_256__81_) );
	INVX1 INVX1_533 ( .A(bloque_in_82_), .Y(_454_) );
	OAI21X1 OAI21X1_676 ( .A(_290__bF_buf11), .B(RAM_entrada_71_bF_buf2), .C(reset_L_bF_buf32), .Y(_455_) );
	AOI21X1 AOI21X1_529 ( .A(_454_), .B(_290__bF_buf10), .C(_455_), .Y(_256__82_) );
	INVX1 INVX1_534 ( .A(bloque_in_83_), .Y(_456_) );
	OAI21X1 OAI21X1_677 ( .A(_290__bF_buf9), .B(RAM_entrada_93_), .C(reset_L_bF_buf31), .Y(_457_) );
	AOI21X1 AOI21X1_530 ( .A(_456_), .B(_290__bF_buf8), .C(_457_), .Y(_256__83_) );
	INVX1 INVX1_535 ( .A(bloque_in_84_), .Y(_458_) );
	OAI21X1 OAI21X1_678 ( .A(_290__bF_buf7), .B(RAM_entrada_89_), .C(reset_L_bF_buf30), .Y(_459_) );
	AOI21X1 AOI21X1_531 ( .A(_458_), .B(_290__bF_buf6), .C(_459_), .Y(_256__84_) );
	INVX1 INVX1_536 ( .A(bloque_in_85_), .Y(_460_) );
	OAI21X1 OAI21X1_679 ( .A(_290__bF_buf5), .B(RAM_entrada_71_bF_buf1), .C(reset_L_bF_buf29), .Y(_461_) );
	AOI21X1 AOI21X1_532 ( .A(_460_), .B(_290__bF_buf4), .C(_461_), .Y(_256__85_) );
	INVX1 INVX1_537 ( .A(bloque_in_86_), .Y(_462_) );
	OAI21X1 OAI21X1_680 ( .A(_290__bF_buf3), .B(RAM_entrada_84_bF_buf1), .C(reset_L_bF_buf28), .Y(_463_) );
	AOI21X1 AOI21X1_533 ( .A(_462_), .B(_290__bF_buf2), .C(_463_), .Y(_256__86_) );
	INVX1 INVX1_538 ( .A(bloque_in_87_), .Y(_464_) );
	OAI21X1 OAI21X1_681 ( .A(_290__bF_buf1), .B(RAM_entrada_85_), .C(reset_L_bF_buf27), .Y(_465_) );
	AOI21X1 AOI21X1_534 ( .A(_464_), .B(_290__bF_buf0), .C(_465_), .Y(_256__87_) );
	INVX1 INVX1_539 ( .A(bloque_in_88_), .Y(_466_) );
	OAI21X1 OAI21X1_682 ( .A(_290__bF_buf15), .B(RAM_entrada_89_), .C(reset_L_bF_buf26), .Y(_467_) );
	AOI21X1 AOI21X1_535 ( .A(_466_), .B(_290__bF_buf14), .C(_467_), .Y(_256__88_) );
	INVX1 INVX1_540 ( .A(bloque_in_89_), .Y(_468_) );
	OAI21X1 OAI21X1_683 ( .A(_290__bF_buf13), .B(RAM_entrada_58_), .C(reset_L_bF_buf25), .Y(_469_) );
	AOI21X1 AOI21X1_536 ( .A(_468_), .B(_290__bF_buf12), .C(_469_), .Y(_256__89_) );
	INVX1 INVX1_541 ( .A(bloque_in_90_), .Y(_470_) );
	OAI21X1 OAI21X1_684 ( .A(_290__bF_buf11), .B(RAM_entrada_58_), .C(reset_L_bF_buf24), .Y(_471_) );
	AOI21X1 AOI21X1_537 ( .A(_470_), .B(_290__bF_buf10), .C(_471_), .Y(_256__90_) );
	INVX1 INVX1_542 ( .A(bloque_in_91_), .Y(_472_) );
	OAI21X1 OAI21X1_685 ( .A(_290__bF_buf9), .B(RAM_entrada_95_), .C(reset_L_bF_buf23), .Y(_473_) );
	AOI21X1 AOI21X1_538 ( .A(_472_), .B(_290__bF_buf8), .C(_473_), .Y(_256__91_) );
	INVX1 INVX1_543 ( .A(bloque_in_92_), .Y(_474_) );
	OAI21X1 OAI21X1_686 ( .A(_290__bF_buf7), .B(RAM_entrada_94_), .C(reset_L_bF_buf22), .Y(_475_) );
	AOI21X1 AOI21X1_539 ( .A(_474_), .B(_290__bF_buf6), .C(_475_), .Y(_256__92_) );
	INVX1 INVX1_544 ( .A(bloque_in_93_), .Y(_476_) );
	OAI21X1 OAI21X1_687 ( .A(_290__bF_buf5), .B(RAM_entrada_71_bF_buf0), .C(reset_L_bF_buf21), .Y(_477_) );
	AOI21X1 AOI21X1_540 ( .A(_476_), .B(_290__bF_buf4), .C(_477_), .Y(_256__93_) );
	INVX1 INVX1_545 ( .A(bloque_in_94_), .Y(_478_) );
	OAI21X1 OAI21X1_688 ( .A(_290__bF_buf3), .B(RAM_entrada_86_), .C(reset_L_bF_buf20), .Y(_479_) );
	AOI21X1 AOI21X1_541 ( .A(_478_), .B(_290__bF_buf2), .C(_479_), .Y(_256__94_) );
	INVX1 INVX1_546 ( .A(bloque_in_95_), .Y(_480_) );
	OAI21X1 OAI21X1_689 ( .A(_290__bF_buf1), .B(RAM_entrada_77_), .C(reset_L_bF_buf19), .Y(_481_) );
	AOI21X1 AOI21X1_542 ( .A(_480_), .B(_290__bF_buf0), .C(_481_), .Y(_256__95_) );
	INVX1 INVX1_547 ( .A(bloque_in_96_), .Y(_482_) );
	OAI21X1 OAI21X1_690 ( .A(_290__bF_buf15), .B(RAM_entrada_88_), .C(reset_L_bF_buf18), .Y(_483_) );
	AOI21X1 AOI21X1_543 ( .A(_482_), .B(_290__bF_buf14), .C(_483_), .Y(_256__96_) );
	INVX1 INVX1_548 ( .A(bloque_in_97_), .Y(_484_) );
	OAI21X1 OAI21X1_691 ( .A(_290__bF_buf13), .B(RAM_entrada_93_), .C(reset_L_bF_buf17), .Y(_485_) );
	AOI21X1 AOI21X1_544 ( .A(_484_), .B(_290__bF_buf12), .C(_485_), .Y(_256__97_) );
	INVX1 INVX1_549 ( .A(bloque_in_98_), .Y(_486_) );
	OAI21X1 OAI21X1_692 ( .A(_290__bF_buf11), .B(RAM_entrada_93_), .C(reset_L_bF_buf16), .Y(_487_) );
	AOI21X1 AOI21X1_545 ( .A(_486_), .B(_290__bF_buf10), .C(_487_), .Y(_256__98_) );
	INVX1 INVX1_550 ( .A(bloque_in_99_), .Y(_488_) );
	OAI21X1 OAI21X1_693 ( .A(_290__bF_buf9), .B(vdd), .C(reset_L_bF_buf15), .Y(_489_) );
	AOI21X1 AOI21X1_546 ( .A(_488_), .B(_290__bF_buf8), .C(_489_), .Y(_256__99_) );
	INVX1 INVX1_551 ( .A(bloque_in_100_), .Y(_490_) );
	OAI21X1 OAI21X1_694 ( .A(_290__bF_buf7), .B(RAM_entrada_89_), .C(reset_L_bF_buf14), .Y(_491_) );
	AOI21X1 AOI21X1_547 ( .A(_490_), .B(_290__bF_buf6), .C(_491_), .Y(_256__100_) );
	INVX1 INVX1_552 ( .A(bloque_in_101_), .Y(_492_) );
	OAI21X1 OAI21X1_695 ( .A(_290__bF_buf5), .B(RAM_entrada_82_), .C(reset_L_bF_buf13), .Y(_493_) );
	AOI21X1 AOI21X1_548 ( .A(_492_), .B(_290__bF_buf4), .C(_493_), .Y(_256__101_) );
	INVX1 INVX1_553 ( .A(bloque_in_102_), .Y(_494_) );
	OAI21X1 OAI21X1_696 ( .A(_290__bF_buf3), .B(RAM_entrada_71_bF_buf3), .C(reset_L_bF_buf12), .Y(_495_) );
	AOI21X1 AOI21X1_549 ( .A(_494_), .B(_290__bF_buf2), .C(_495_), .Y(_256__102_) );
	INVX1 INVX1_554 ( .A(bloque_in_103_), .Y(_496_) );
	OAI21X1 OAI21X1_697 ( .A(_290__bF_buf1), .B(RAM_entrada_71_bF_buf2), .C(reset_L_bF_buf11), .Y(_497_) );
	AOI21X1 AOI21X1_550 ( .A(_496_), .B(_290__bF_buf0), .C(_497_), .Y(_256__103_) );
	INVX1 INVX1_555 ( .A(bloque_in_104_), .Y(_498_) );
	OAI21X1 OAI21X1_698 ( .A(_290__bF_buf15), .B(RAM_entrada_92_), .C(reset_L_bF_buf10), .Y(_499_) );
	AOI21X1 AOI21X1_551 ( .A(_498_), .B(_290__bF_buf14), .C(_499_), .Y(_256__104_) );
	INVX1 INVX1_556 ( .A(bloque_in_105_), .Y(_500_) );
	OAI21X1 OAI21X1_699 ( .A(_290__bF_buf13), .B(RAM_entrada_88_), .C(reset_L_bF_buf9), .Y(_501_) );
	AOI21X1 AOI21X1_552 ( .A(_500_), .B(_290__bF_buf12), .C(_501_), .Y(_256__105_) );
	INVX1 INVX1_557 ( .A(bloque_in_106_), .Y(_502_) );
	OAI21X1 OAI21X1_700 ( .A(_290__bF_buf11), .B(RAM_entrada_88_), .C(reset_L_bF_buf8), .Y(_503_) );
	AOI21X1 AOI21X1_553 ( .A(_502_), .B(_290__bF_buf10), .C(_503_), .Y(_256__106_) );
	INVX1 INVX1_558 ( .A(bloque_in_107_), .Y(_504_) );
	OAI21X1 OAI21X1_701 ( .A(_290__bF_buf9), .B(vdd), .C(reset_L_bF_buf7), .Y(_505_) );
	AOI21X1 AOI21X1_554 ( .A(_504_), .B(_290__bF_buf8), .C(_505_), .Y(_256__107_) );
	INVX1 INVX1_559 ( .A(bloque_in_108_), .Y(_506_) );
	OAI21X1 OAI21X1_702 ( .A(_290__bF_buf7), .B(RAM_entrada_84_bF_buf0), .C(reset_L_bF_buf6), .Y(_507_) );
	AOI21X1 AOI21X1_555 ( .A(_506_), .B(_290__bF_buf6), .C(_507_), .Y(_256__108_) );
	INVX1 INVX1_560 ( .A(bloque_in_109_), .Y(_508_) );
	OAI21X1 OAI21X1_703 ( .A(_290__bF_buf5), .B(RAM_entrada_77_), .C(reset_L_bF_buf5), .Y(_509_) );
	AOI21X1 AOI21X1_556 ( .A(_508_), .B(_290__bF_buf4), .C(_509_), .Y(_256__109_) );
	INVX1 INVX1_561 ( .A(bloque_in_110_), .Y(_510_) );
	OAI21X1 OAI21X1_704 ( .A(_290__bF_buf3), .B(RAM_entrada_89_), .C(reset_L_bF_buf4), .Y(_511_) );
	AOI21X1 AOI21X1_557 ( .A(_510_), .B(_290__bF_buf2), .C(_511_), .Y(_256__110_) );
	INVX1 INVX1_562 ( .A(bloque_in_111_), .Y(_512_) );
	OAI21X1 OAI21X1_705 ( .A(_290__bF_buf1), .B(RAM_entrada_88_), .C(reset_L_bF_buf3), .Y(_513_) );
	AOI21X1 AOI21X1_558 ( .A(_512_), .B(_290__bF_buf0), .C(_513_), .Y(_256__111_) );
	INVX1 INVX1_563 ( .A(bloque_in_112_), .Y(_514_) );
	OAI21X1 OAI21X1_706 ( .A(_290__bF_buf15), .B(RAM_entrada_85_), .C(reset_L_bF_buf2), .Y(_515_) );
	AOI21X1 AOI21X1_559 ( .A(_514_), .B(_290__bF_buf14), .C(_515_), .Y(_256__112_) );
	INVX1 INVX1_564 ( .A(bloque_in_113_), .Y(_516_) );
	OAI21X1 OAI21X1_707 ( .A(_290__bF_buf13), .B(RAM_entrada_89_), .C(reset_L_bF_buf1), .Y(_517_) );
	AOI21X1 AOI21X1_560 ( .A(_516_), .B(_290__bF_buf12), .C(_517_), .Y(_256__113_) );
	INVX1 INVX1_565 ( .A(bloque_in_114_), .Y(_518_) );
	OAI21X1 OAI21X1_708 ( .A(_290__bF_buf11), .B(RAM_entrada_82_), .C(reset_L_bF_buf0), .Y(_519_) );
	AOI21X1 AOI21X1_561 ( .A(_518_), .B(_290__bF_buf10), .C(_519_), .Y(_256__114_) );
	INVX1 INVX1_566 ( .A(bloque_in_115_), .Y(_520_) );
	OAI21X1 OAI21X1_709 ( .A(_290__bF_buf9), .B(RAM_entrada_84_bF_buf3), .C(reset_L_bF_buf49), .Y(_521_) );
	AOI21X1 AOI21X1_562 ( .A(_520_), .B(_290__bF_buf8), .C(_521_), .Y(_256__115_) );
	INVX1 INVX1_567 ( .A(bloque_in_116_), .Y(_522_) );
	OAI21X1 OAI21X1_710 ( .A(_290__bF_buf7), .B(RAM_entrada_84_bF_buf2), .C(reset_L_bF_buf48), .Y(_523_) );
	AOI21X1 AOI21X1_563 ( .A(_522_), .B(_290__bF_buf6), .C(_523_), .Y(_256__116_) );
	INVX1 INVX1_568 ( .A(bloque_in_117_), .Y(_524_) );
	OAI21X1 OAI21X1_711 ( .A(_290__bF_buf5), .B(RAM_entrada_85_), .C(reset_L_bF_buf47), .Y(_525_) );
	AOI21X1 AOI21X1_564 ( .A(_524_), .B(_290__bF_buf4), .C(_525_), .Y(_256__117_) );
	INVX1 INVX1_569 ( .A(bloque_in_118_), .Y(_526_) );
	OAI21X1 OAI21X1_712 ( .A(_290__bF_buf3), .B(RAM_entrada_86_), .C(reset_L_bF_buf46), .Y(_527_) );
	AOI21X1 AOI21X1_565 ( .A(_526_), .B(_290__bF_buf2), .C(_527_), .Y(_256__118_) );
	INVX1 INVX1_570 ( .A(bloque_in_119_), .Y(_528_) );
	OAI21X1 OAI21X1_713 ( .A(_290__bF_buf1), .B(gnd), .C(reset_L_bF_buf45), .Y(_529_) );
	AOI21X1 AOI21X1_566 ( .A(_528_), .B(_290__bF_buf0), .C(_529_), .Y(_256__119_) );
	INVX1 INVX1_571 ( .A(bloque_in_120_), .Y(_530_) );
	OAI21X1 OAI21X1_714 ( .A(_290__bF_buf15), .B(RAM_entrada_88_), .C(reset_L_bF_buf44), .Y(_531_) );
	AOI21X1 AOI21X1_567 ( .A(_530_), .B(_290__bF_buf14), .C(_531_), .Y(_256__120_) );
	INVX1 INVX1_572 ( .A(bloque_in_121_), .Y(_532_) );
	OAI21X1 OAI21X1_715 ( .A(_290__bF_buf13), .B(RAM_entrada_89_), .C(reset_L_bF_buf43), .Y(_533_) );
	AOI21X1 AOI21X1_568 ( .A(_532_), .B(_290__bF_buf12), .C(_533_), .Y(_256__121_) );
	INVX1 INVX1_573 ( .A(bloque_in_122_), .Y(_534_) );
	OAI21X1 OAI21X1_716 ( .A(_290__bF_buf11), .B(RAM_entrada_94_), .C(reset_L_bF_buf42), .Y(_535_) );
	AOI21X1 AOI21X1_569 ( .A(_534_), .B(_290__bF_buf10), .C(_535_), .Y(_256__122_) );
	INVX1 INVX1_574 ( .A(bloque_in_123_), .Y(_536_) );
	OAI21X1 OAI21X1_717 ( .A(_290__bF_buf9), .B(vdd), .C(reset_L_bF_buf41), .Y(_537_) );
	AOI21X1 AOI21X1_570 ( .A(_536_), .B(_290__bF_buf8), .C(_537_), .Y(_256__123_) );
	INVX1 INVX1_575 ( .A(bloque_in_124_), .Y(_538_) );
	OAI21X1 OAI21X1_718 ( .A(_290__bF_buf7), .B(RAM_entrada_92_), .C(reset_L_bF_buf40), .Y(_539_) );
	AOI21X1 AOI21X1_571 ( .A(_538_), .B(_290__bF_buf6), .C(_539_), .Y(_256__124_) );
	INVX1 INVX1_576 ( .A(bloque_in_125_), .Y(_540_) );
	OAI21X1 OAI21X1_719 ( .A(_290__bF_buf5), .B(RAM_entrada_93_), .C(reset_L_bF_buf39), .Y(_541_) );
	AOI21X1 AOI21X1_572 ( .A(_540_), .B(_290__bF_buf4), .C(_541_), .Y(_256__125_) );
	INVX1 INVX1_577 ( .A(bloque_in_126_), .Y(_542_) );
	OAI21X1 OAI21X1_720 ( .A(_290__bF_buf3), .B(RAM_entrada_94_), .C(reset_L_bF_buf38), .Y(_543_) );
	AOI21X1 AOI21X1_573 ( .A(_542_), .B(_290__bF_buf2), .C(_543_), .Y(_256__126_) );
	INVX1 INVX1_578 ( .A(bloque_in_127_), .Y(_544_) );
	OAI21X1 OAI21X1_721 ( .A(_290__bF_buf1), .B(RAM_entrada_95_), .C(reset_L_bF_buf37), .Y(_545_) );
	AOI21X1 AOI21X1_574 ( .A(_544_), .B(_290__bF_buf0), .C(_545_), .Y(_256__127_) );
	DFFPOSX1 DFFPOSX1_541 ( .CLK(clk_bF_buf29), .D(_256__0_), .Q(bloque_in_0_) );
	DFFPOSX1 DFFPOSX1_542 ( .CLK(clk_bF_buf28), .D(_256__1_), .Q(bloque_in_1_) );
	DFFPOSX1 DFFPOSX1_543 ( .CLK(clk_bF_buf27), .D(_256__2_), .Q(bloque_in_2_) );
	DFFPOSX1 DFFPOSX1_544 ( .CLK(clk_bF_buf26), .D(_256__3_), .Q(bloque_in_3_) );
	DFFPOSX1 DFFPOSX1_545 ( .CLK(clk_bF_buf25), .D(_256__4_), .Q(bloque_in_4_) );
	DFFPOSX1 DFFPOSX1_546 ( .CLK(clk_bF_buf24), .D(_256__5_), .Q(bloque_in_5_) );
	DFFPOSX1 DFFPOSX1_547 ( .CLK(clk_bF_buf23), .D(_256__6_), .Q(bloque_in_6_) );
	DFFPOSX1 DFFPOSX1_548 ( .CLK(clk_bF_buf22), .D(_256__7_), .Q(bloque_in_7_) );
	DFFPOSX1 DFFPOSX1_549 ( .CLK(clk_bF_buf21), .D(_256__8_), .Q(bloque_in_8_) );
	DFFPOSX1 DFFPOSX1_550 ( .CLK(clk_bF_buf20), .D(_256__9_), .Q(bloque_in_9_) );
	DFFPOSX1 DFFPOSX1_551 ( .CLK(clk_bF_buf19), .D(_256__10_), .Q(bloque_in_10_) );
	DFFPOSX1 DFFPOSX1_552 ( .CLK(clk_bF_buf18), .D(_256__11_), .Q(bloque_in_11_) );
	DFFPOSX1 DFFPOSX1_553 ( .CLK(clk_bF_buf17), .D(_256__12_), .Q(bloque_in_12_) );
	DFFPOSX1 DFFPOSX1_554 ( .CLK(clk_bF_buf16), .D(_256__13_), .Q(bloque_in_13_) );
	DFFPOSX1 DFFPOSX1_555 ( .CLK(clk_bF_buf15), .D(_256__14_), .Q(bloque_in_14_) );
	DFFPOSX1 DFFPOSX1_556 ( .CLK(clk_bF_buf14), .D(_256__15_), .Q(bloque_in_15_) );
	DFFPOSX1 DFFPOSX1_557 ( .CLK(clk_bF_buf13), .D(_256__16_), .Q(bloque_in_16_) );
	DFFPOSX1 DFFPOSX1_558 ( .CLK(clk_bF_buf12), .D(_256__17_), .Q(bloque_in_17_) );
	DFFPOSX1 DFFPOSX1_559 ( .CLK(clk_bF_buf11), .D(_256__18_), .Q(bloque_in_18_) );
	DFFPOSX1 DFFPOSX1_560 ( .CLK(clk_bF_buf10), .D(_256__19_), .Q(bloque_in_19_) );
	DFFPOSX1 DFFPOSX1_561 ( .CLK(clk_bF_buf9), .D(_256__20_), .Q(bloque_in_20_) );
	DFFPOSX1 DFFPOSX1_562 ( .CLK(clk_bF_buf8), .D(_256__21_), .Q(bloque_in_21_) );
	DFFPOSX1 DFFPOSX1_563 ( .CLK(clk_bF_buf7), .D(_256__22_), .Q(bloque_in_22_) );
	DFFPOSX1 DFFPOSX1_564 ( .CLK(clk_bF_buf6), .D(_256__23_), .Q(bloque_in_23_) );
	DFFPOSX1 DFFPOSX1_565 ( .CLK(clk_bF_buf5), .D(_256__24_), .Q(bloque_in_24_) );
	DFFPOSX1 DFFPOSX1_566 ( .CLK(clk_bF_buf4), .D(_256__25_), .Q(bloque_in_25_) );
	DFFPOSX1 DFFPOSX1_567 ( .CLK(clk_bF_buf3), .D(_256__26_), .Q(bloque_in_26_) );
	DFFPOSX1 DFFPOSX1_568 ( .CLK(clk_bF_buf2), .D(_256__27_), .Q(bloque_in_27_) );
	DFFPOSX1 DFFPOSX1_569 ( .CLK(clk_bF_buf1), .D(_256__28_), .Q(bloque_in_28_) );
	DFFPOSX1 DFFPOSX1_570 ( .CLK(clk_bF_buf0), .D(_256__29_), .Q(bloque_in_29_) );
	DFFPOSX1 DFFPOSX1_571 ( .CLK(clk_bF_buf113), .D(_256__30_), .Q(bloque_in_30_) );
	DFFPOSX1 DFFPOSX1_572 ( .CLK(clk_bF_buf112), .D(_256__31_), .Q(bloque_in_31_) );
	DFFPOSX1 DFFPOSX1_573 ( .CLK(clk_bF_buf111), .D(_256__32_), .Q(bloque_in_32_) );
	DFFPOSX1 DFFPOSX1_574 ( .CLK(clk_bF_buf110), .D(_256__33_), .Q(bloque_in_33_) );
	DFFPOSX1 DFFPOSX1_575 ( .CLK(clk_bF_buf109), .D(_256__34_), .Q(bloque_in_34_) );
	DFFPOSX1 DFFPOSX1_576 ( .CLK(clk_bF_buf108), .D(_256__35_), .Q(bloque_in_35_) );
	DFFPOSX1 DFFPOSX1_577 ( .CLK(clk_bF_buf107), .D(_256__36_), .Q(bloque_in_36_) );
	DFFPOSX1 DFFPOSX1_578 ( .CLK(clk_bF_buf106), .D(_256__37_), .Q(bloque_in_37_) );
	DFFPOSX1 DFFPOSX1_579 ( .CLK(clk_bF_buf105), .D(_256__38_), .Q(bloque_in_38_) );
	DFFPOSX1 DFFPOSX1_580 ( .CLK(clk_bF_buf104), .D(_256__39_), .Q(bloque_in_39_) );
	DFFPOSX1 DFFPOSX1_581 ( .CLK(clk_bF_buf103), .D(_256__40_), .Q(bloque_in_40_) );
	DFFPOSX1 DFFPOSX1_582 ( .CLK(clk_bF_buf102), .D(_256__41_), .Q(bloque_in_41_) );
	DFFPOSX1 DFFPOSX1_583 ( .CLK(clk_bF_buf101), .D(_256__42_), .Q(bloque_in_42_) );
	DFFPOSX1 DFFPOSX1_584 ( .CLK(clk_bF_buf100), .D(_256__43_), .Q(bloque_in_43_) );
	DFFPOSX1 DFFPOSX1_585 ( .CLK(clk_bF_buf99), .D(_256__44_), .Q(bloque_in_44_) );
	DFFPOSX1 DFFPOSX1_586 ( .CLK(clk_bF_buf98), .D(_256__45_), .Q(bloque_in_45_) );
	DFFPOSX1 DFFPOSX1_587 ( .CLK(clk_bF_buf97), .D(_256__46_), .Q(bloque_in_46_) );
	DFFPOSX1 DFFPOSX1_588 ( .CLK(clk_bF_buf96), .D(_256__47_), .Q(bloque_in_47_) );
	DFFPOSX1 DFFPOSX1_589 ( .CLK(clk_bF_buf95), .D(_256__48_), .Q(bloque_in_48_) );
	DFFPOSX1 DFFPOSX1_590 ( .CLK(clk_bF_buf94), .D(_256__49_), .Q(bloque_in_49_) );
	DFFPOSX1 DFFPOSX1_591 ( .CLK(clk_bF_buf93), .D(_256__50_), .Q(bloque_in_50_) );
	DFFPOSX1 DFFPOSX1_592 ( .CLK(clk_bF_buf92), .D(_256__51_), .Q(bloque_in_51_) );
	DFFPOSX1 DFFPOSX1_593 ( .CLK(clk_bF_buf91), .D(_256__52_), .Q(bloque_in_52_) );
	DFFPOSX1 DFFPOSX1_594 ( .CLK(clk_bF_buf90), .D(_256__53_), .Q(bloque_in_53_) );
	DFFPOSX1 DFFPOSX1_595 ( .CLK(clk_bF_buf89), .D(_256__54_), .Q(bloque_in_54_) );
	DFFPOSX1 DFFPOSX1_596 ( .CLK(clk_bF_buf88), .D(_256__55_), .Q(bloque_in_55_) );
	DFFPOSX1 DFFPOSX1_597 ( .CLK(clk_bF_buf87), .D(_256__56_), .Q(bloque_in_56_) );
	DFFPOSX1 DFFPOSX1_598 ( .CLK(clk_bF_buf86), .D(_256__57_), .Q(bloque_in_57_) );
	DFFPOSX1 DFFPOSX1_599 ( .CLK(clk_bF_buf85), .D(_256__58_), .Q(bloque_in_58_) );
	DFFPOSX1 DFFPOSX1_600 ( .CLK(clk_bF_buf84), .D(_256__59_), .Q(bloque_in_59_) );
	DFFPOSX1 DFFPOSX1_601 ( .CLK(clk_bF_buf83), .D(_256__60_), .Q(bloque_in_60_) );
	DFFPOSX1 DFFPOSX1_602 ( .CLK(clk_bF_buf82), .D(_256__61_), .Q(bloque_in_61_) );
	DFFPOSX1 DFFPOSX1_603 ( .CLK(clk_bF_buf81), .D(_256__62_), .Q(bloque_in_62_) );
	DFFPOSX1 DFFPOSX1_604 ( .CLK(clk_bF_buf80), .D(_256__63_), .Q(bloque_in_63_) );
	DFFPOSX1 DFFPOSX1_605 ( .CLK(clk_bF_buf79), .D(_256__64_), .Q(bloque_in_64_) );
	DFFPOSX1 DFFPOSX1_606 ( .CLK(clk_bF_buf78), .D(_256__65_), .Q(bloque_in_65_) );
	DFFPOSX1 DFFPOSX1_607 ( .CLK(clk_bF_buf77), .D(_256__66_), .Q(bloque_in_66_) );
	DFFPOSX1 DFFPOSX1_608 ( .CLK(clk_bF_buf76), .D(_256__67_), .Q(bloque_in_67_) );
	DFFPOSX1 DFFPOSX1_609 ( .CLK(clk_bF_buf75), .D(_256__68_), .Q(bloque_in_68_) );
	DFFPOSX1 DFFPOSX1_610 ( .CLK(clk_bF_buf74), .D(_256__69_), .Q(bloque_in_69_) );
	DFFPOSX1 DFFPOSX1_611 ( .CLK(clk_bF_buf73), .D(_256__70_), .Q(bloque_in_70_) );
	DFFPOSX1 DFFPOSX1_612 ( .CLK(clk_bF_buf72), .D(_256__71_), .Q(bloque_in_71_) );
	DFFPOSX1 DFFPOSX1_613 ( .CLK(clk_bF_buf71), .D(_256__72_), .Q(bloque_in_72_) );
	DFFPOSX1 DFFPOSX1_614 ( .CLK(clk_bF_buf70), .D(_256__73_), .Q(bloque_in_73_) );
	DFFPOSX1 DFFPOSX1_615 ( .CLK(clk_bF_buf69), .D(_256__74_), .Q(bloque_in_74_) );
	DFFPOSX1 DFFPOSX1_616 ( .CLK(clk_bF_buf68), .D(_256__75_), .Q(bloque_in_75_) );
	DFFPOSX1 DFFPOSX1_617 ( .CLK(clk_bF_buf67), .D(_256__76_), .Q(bloque_in_76_) );
	DFFPOSX1 DFFPOSX1_618 ( .CLK(clk_bF_buf66), .D(_256__77_), .Q(bloque_in_77_) );
	DFFPOSX1 DFFPOSX1_619 ( .CLK(clk_bF_buf65), .D(_256__78_), .Q(bloque_in_78_) );
	DFFPOSX1 DFFPOSX1_620 ( .CLK(clk_bF_buf64), .D(_256__79_), .Q(bloque_in_79_) );
	DFFPOSX1 DFFPOSX1_621 ( .CLK(clk_bF_buf63), .D(_256__80_), .Q(bloque_in_80_) );
	DFFPOSX1 DFFPOSX1_622 ( .CLK(clk_bF_buf62), .D(_256__81_), .Q(bloque_in_81_) );
	DFFPOSX1 DFFPOSX1_623 ( .CLK(clk_bF_buf61), .D(_256__82_), .Q(bloque_in_82_) );
	DFFPOSX1 DFFPOSX1_624 ( .CLK(clk_bF_buf60), .D(_256__83_), .Q(bloque_in_83_) );
	DFFPOSX1 DFFPOSX1_625 ( .CLK(clk_bF_buf59), .D(_256__84_), .Q(bloque_in_84_) );
	DFFPOSX1 DFFPOSX1_626 ( .CLK(clk_bF_buf58), .D(_256__85_), .Q(bloque_in_85_) );
	DFFPOSX1 DFFPOSX1_627 ( .CLK(clk_bF_buf57), .D(_256__86_), .Q(bloque_in_86_) );
	DFFPOSX1 DFFPOSX1_628 ( .CLK(clk_bF_buf56), .D(_256__87_), .Q(bloque_in_87_) );
	DFFPOSX1 DFFPOSX1_629 ( .CLK(clk_bF_buf55), .D(_256__88_), .Q(bloque_in_88_) );
	DFFPOSX1 DFFPOSX1_630 ( .CLK(clk_bF_buf54), .D(_256__89_), .Q(bloque_in_89_) );
	DFFPOSX1 DFFPOSX1_631 ( .CLK(clk_bF_buf53), .D(_256__90_), .Q(bloque_in_90_) );
	DFFPOSX1 DFFPOSX1_632 ( .CLK(clk_bF_buf52), .D(_256__91_), .Q(bloque_in_91_) );
	DFFPOSX1 DFFPOSX1_633 ( .CLK(clk_bF_buf51), .D(_256__92_), .Q(bloque_in_92_) );
	DFFPOSX1 DFFPOSX1_634 ( .CLK(clk_bF_buf50), .D(_256__93_), .Q(bloque_in_93_) );
	DFFPOSX1 DFFPOSX1_635 ( .CLK(clk_bF_buf49), .D(_256__94_), .Q(bloque_in_94_) );
	DFFPOSX1 DFFPOSX1_636 ( .CLK(clk_bF_buf48), .D(_256__95_), .Q(bloque_in_95_) );
	DFFPOSX1 DFFPOSX1_637 ( .CLK(clk_bF_buf47), .D(_256__96_), .Q(bloque_in_96_) );
	DFFPOSX1 DFFPOSX1_638 ( .CLK(clk_bF_buf46), .D(_256__97_), .Q(bloque_in_97_) );
	DFFPOSX1 DFFPOSX1_639 ( .CLK(clk_bF_buf45), .D(_256__98_), .Q(bloque_in_98_) );
	DFFPOSX1 DFFPOSX1_640 ( .CLK(clk_bF_buf44), .D(_256__99_), .Q(bloque_in_99_) );
	DFFPOSX1 DFFPOSX1_641 ( .CLK(clk_bF_buf43), .D(_256__100_), .Q(bloque_in_100_) );
	DFFPOSX1 DFFPOSX1_642 ( .CLK(clk_bF_buf42), .D(_256__101_), .Q(bloque_in_101_) );
	DFFPOSX1 DFFPOSX1_643 ( .CLK(clk_bF_buf41), .D(_256__102_), .Q(bloque_in_102_) );
	DFFPOSX1 DFFPOSX1_644 ( .CLK(clk_bF_buf40), .D(_256__103_), .Q(bloque_in_103_) );
	DFFPOSX1 DFFPOSX1_645 ( .CLK(clk_bF_buf39), .D(_256__104_), .Q(bloque_in_104_) );
	DFFPOSX1 DFFPOSX1_646 ( .CLK(clk_bF_buf38), .D(_256__105_), .Q(bloque_in_105_) );
	DFFPOSX1 DFFPOSX1_647 ( .CLK(clk_bF_buf37), .D(_256__106_), .Q(bloque_in_106_) );
	DFFPOSX1 DFFPOSX1_648 ( .CLK(clk_bF_buf36), .D(_256__107_), .Q(bloque_in_107_) );
	DFFPOSX1 DFFPOSX1_649 ( .CLK(clk_bF_buf35), .D(_256__108_), .Q(bloque_in_108_) );
	DFFPOSX1 DFFPOSX1_650 ( .CLK(clk_bF_buf34), .D(_256__109_), .Q(bloque_in_109_) );
	DFFPOSX1 DFFPOSX1_651 ( .CLK(clk_bF_buf33), .D(_256__110_), .Q(bloque_in_110_) );
	DFFPOSX1 DFFPOSX1_652 ( .CLK(clk_bF_buf32), .D(_256__111_), .Q(bloque_in_111_) );
	DFFPOSX1 DFFPOSX1_653 ( .CLK(clk_bF_buf31), .D(_256__112_), .Q(bloque_in_112_) );
	DFFPOSX1 DFFPOSX1_654 ( .CLK(clk_bF_buf30), .D(_256__113_), .Q(bloque_in_113_) );
	DFFPOSX1 DFFPOSX1_655 ( .CLK(clk_bF_buf29), .D(_256__114_), .Q(bloque_in_114_) );
	DFFPOSX1 DFFPOSX1_656 ( .CLK(clk_bF_buf28), .D(_256__115_), .Q(bloque_in_115_) );
	DFFPOSX1 DFFPOSX1_657 ( .CLK(clk_bF_buf27), .D(_256__116_), .Q(bloque_in_116_) );
	DFFPOSX1 DFFPOSX1_658 ( .CLK(clk_bF_buf26), .D(_256__117_), .Q(bloque_in_117_) );
	DFFPOSX1 DFFPOSX1_659 ( .CLK(clk_bF_buf25), .D(_256__118_), .Q(bloque_in_118_) );
	DFFPOSX1 DFFPOSX1_660 ( .CLK(clk_bF_buf24), .D(_256__119_), .Q(bloque_in_119_) );
	DFFPOSX1 DFFPOSX1_661 ( .CLK(clk_bF_buf23), .D(_256__120_), .Q(bloque_in_120_) );
	DFFPOSX1 DFFPOSX1_662 ( .CLK(clk_bF_buf22), .D(_256__121_), .Q(bloque_in_121_) );
	DFFPOSX1 DFFPOSX1_663 ( .CLK(clk_bF_buf21), .D(_256__122_), .Q(bloque_in_122_) );
	DFFPOSX1 DFFPOSX1_664 ( .CLK(clk_bF_buf20), .D(_256__123_), .Q(bloque_in_123_) );
	DFFPOSX1 DFFPOSX1_665 ( .CLK(clk_bF_buf19), .D(_256__124_), .Q(bloque_in_124_) );
	DFFPOSX1 DFFPOSX1_666 ( .CLK(clk_bF_buf18), .D(_256__125_), .Q(bloque_in_125_) );
	DFFPOSX1 DFFPOSX1_667 ( .CLK(clk_bF_buf17), .D(_256__126_), .Q(bloque_in_126_) );
	DFFPOSX1 DFFPOSX1_668 ( .CLK(clk_bF_buf16), .D(_256__127_), .Q(bloque_in_127_) );
	DFFPOSX1 DFFPOSX1_669 ( .CLK(clk_bF_buf15), .D(_257__0_), .Q(bloque_in_1_0_) );
	DFFPOSX1 DFFPOSX1_670 ( .CLK(clk_bF_buf14), .D(_257__1_), .Q(bloque_in_1_1_) );
	DFFPOSX1 DFFPOSX1_671 ( .CLK(clk_bF_buf13), .D(_257__2_), .Q(bloque_in_1_2_) );
	DFFPOSX1 DFFPOSX1_672 ( .CLK(clk_bF_buf12), .D(_257__3_), .Q(bloque_in_1_3_) );
	DFFPOSX1 DFFPOSX1_673 ( .CLK(clk_bF_buf11), .D(_257__4_), .Q(bloque_in_1_4_) );
	DFFPOSX1 DFFPOSX1_674 ( .CLK(clk_bF_buf10), .D(_257__5_), .Q(bloque_in_1_5_) );
	DFFPOSX1 DFFPOSX1_675 ( .CLK(clk_bF_buf9), .D(_257__6_), .Q(bloque_in_1_6_) );
	DFFPOSX1 DFFPOSX1_676 ( .CLK(clk_bF_buf8), .D(_257__7_), .Q(bloque_in_1_7_) );
	DFFPOSX1 DFFPOSX1_677 ( .CLK(clk_bF_buf7), .D(_257__8_), .Q(bloque_in_1_8_) );
	DFFPOSX1 DFFPOSX1_678 ( .CLK(clk_bF_buf6), .D(_257__9_), .Q(bloque_in_1_9_) );
	DFFPOSX1 DFFPOSX1_679 ( .CLK(clk_bF_buf5), .D(_257__10_), .Q(bloque_in_1_10_) );
	DFFPOSX1 DFFPOSX1_680 ( .CLK(clk_bF_buf4), .D(_257__11_), .Q(bloque_in_1_11_) );
	DFFPOSX1 DFFPOSX1_681 ( .CLK(clk_bF_buf3), .D(_257__12_), .Q(bloque_in_1_12_) );
	DFFPOSX1 DFFPOSX1_682 ( .CLK(clk_bF_buf2), .D(_257__13_), .Q(bloque_in_1_13_) );
	DFFPOSX1 DFFPOSX1_683 ( .CLK(clk_bF_buf1), .D(_257__14_), .Q(bloque_in_1_14_) );
	DFFPOSX1 DFFPOSX1_684 ( .CLK(clk_bF_buf0), .D(_257__15_), .Q(bloque_in_1_15_) );
	DFFPOSX1 DFFPOSX1_685 ( .CLK(clk_bF_buf113), .D(_257__16_), .Q(bloque_in_1_16_) );
	DFFPOSX1 DFFPOSX1_686 ( .CLK(clk_bF_buf112), .D(_257__17_), .Q(bloque_in_1_17_) );
	DFFPOSX1 DFFPOSX1_687 ( .CLK(clk_bF_buf111), .D(_257__18_), .Q(bloque_in_1_18_) );
	DFFPOSX1 DFFPOSX1_688 ( .CLK(clk_bF_buf110), .D(_257__19_), .Q(bloque_in_1_19_) );
	DFFPOSX1 DFFPOSX1_689 ( .CLK(clk_bF_buf109), .D(_257__20_), .Q(bloque_in_1_20_) );
	DFFPOSX1 DFFPOSX1_690 ( .CLK(clk_bF_buf108), .D(_257__21_), .Q(bloque_in_1_21_) );
	DFFPOSX1 DFFPOSX1_691 ( .CLK(clk_bF_buf107), .D(_257__22_), .Q(bloque_in_1_22_) );
	DFFPOSX1 DFFPOSX1_692 ( .CLK(clk_bF_buf106), .D(_257__23_), .Q(bloque_in_1_23_) );
	DFFPOSX1 DFFPOSX1_693 ( .CLK(clk_bF_buf105), .D(_257__24_), .Q(bloque_in_1_24_) );
	DFFPOSX1 DFFPOSX1_694 ( .CLK(clk_bF_buf104), .D(_257__25_), .Q(bloque_in_1_25_) );
	DFFPOSX1 DFFPOSX1_695 ( .CLK(clk_bF_buf103), .D(_257__26_), .Q(bloque_in_1_26_) );
	DFFPOSX1 DFFPOSX1_696 ( .CLK(clk_bF_buf102), .D(_257__27_), .Q(bloque_in_1_27_) );
	DFFPOSX1 DFFPOSX1_697 ( .CLK(clk_bF_buf101), .D(_257__28_), .Q(bloque_in_1_28_) );
	DFFPOSX1 DFFPOSX1_698 ( .CLK(clk_bF_buf100), .D(_257__29_), .Q(bloque_in_1_29_) );
	DFFPOSX1 DFFPOSX1_699 ( .CLK(clk_bF_buf99), .D(_257__30_), .Q(bloque_in_1_30_) );
	DFFPOSX1 DFFPOSX1_700 ( .CLK(clk_bF_buf98), .D(_257__31_), .Q(bloque_in_1_31_) );
	DFFPOSX1 DFFPOSX1_701 ( .CLK(clk_bF_buf97), .D(_257__32_), .Q(bloque_in_1_32_) );
	DFFPOSX1 DFFPOSX1_702 ( .CLK(clk_bF_buf96), .D(_257__33_), .Q(bloque_in_1_33_) );
	DFFPOSX1 DFFPOSX1_703 ( .CLK(clk_bF_buf95), .D(_257__34_), .Q(bloque_in_1_34_) );
	DFFPOSX1 DFFPOSX1_704 ( .CLK(clk_bF_buf94), .D(_257__35_), .Q(bloque_in_1_35_) );
	DFFPOSX1 DFFPOSX1_705 ( .CLK(clk_bF_buf93), .D(_257__36_), .Q(bloque_in_1_36_) );
	DFFPOSX1 DFFPOSX1_706 ( .CLK(clk_bF_buf92), .D(_257__37_), .Q(bloque_in_1_37_) );
	DFFPOSX1 DFFPOSX1_707 ( .CLK(clk_bF_buf91), .D(_257__38_), .Q(bloque_in_1_38_) );
	DFFPOSX1 DFFPOSX1_708 ( .CLK(clk_bF_buf90), .D(_257__39_), .Q(bloque_in_1_39_) );
	DFFPOSX1 DFFPOSX1_709 ( .CLK(clk_bF_buf89), .D(_257__40_), .Q(bloque_in_1_40_) );
	DFFPOSX1 DFFPOSX1_710 ( .CLK(clk_bF_buf88), .D(_257__41_), .Q(bloque_in_1_41_) );
	DFFPOSX1 DFFPOSX1_711 ( .CLK(clk_bF_buf87), .D(_257__42_), .Q(bloque_in_1_42_) );
	DFFPOSX1 DFFPOSX1_712 ( .CLK(clk_bF_buf86), .D(_257__43_), .Q(bloque_in_1_43_) );
	DFFPOSX1 DFFPOSX1_713 ( .CLK(clk_bF_buf85), .D(_257__44_), .Q(bloque_in_1_44_) );
	DFFPOSX1 DFFPOSX1_714 ( .CLK(clk_bF_buf84), .D(_257__45_), .Q(bloque_in_1_45_) );
	DFFPOSX1 DFFPOSX1_715 ( .CLK(clk_bF_buf83), .D(_257__46_), .Q(bloque_in_1_46_) );
	DFFPOSX1 DFFPOSX1_716 ( .CLK(clk_bF_buf82), .D(_257__47_), .Q(bloque_in_1_47_) );
	DFFPOSX1 DFFPOSX1_717 ( .CLK(clk_bF_buf81), .D(_257__48_), .Q(bloque_in_1_48_) );
	DFFPOSX1 DFFPOSX1_718 ( .CLK(clk_bF_buf80), .D(_257__49_), .Q(bloque_in_1_49_) );
	DFFPOSX1 DFFPOSX1_719 ( .CLK(clk_bF_buf79), .D(_257__50_), .Q(bloque_in_1_50_) );
	DFFPOSX1 DFFPOSX1_720 ( .CLK(clk_bF_buf78), .D(_257__51_), .Q(bloque_in_1_51_) );
	DFFPOSX1 DFFPOSX1_721 ( .CLK(clk_bF_buf77), .D(_257__52_), .Q(bloque_in_1_52_) );
	DFFPOSX1 DFFPOSX1_722 ( .CLK(clk_bF_buf76), .D(_257__53_), .Q(bloque_in_1_53_) );
	DFFPOSX1 DFFPOSX1_723 ( .CLK(clk_bF_buf75), .D(_257__54_), .Q(bloque_in_1_54_) );
	DFFPOSX1 DFFPOSX1_724 ( .CLK(clk_bF_buf74), .D(_257__55_), .Q(bloque_in_1_55_) );
	DFFPOSX1 DFFPOSX1_725 ( .CLK(clk_bF_buf73), .D(_257__56_), .Q(bloque_in_1_56_) );
	DFFPOSX1 DFFPOSX1_726 ( .CLK(clk_bF_buf72), .D(_257__57_), .Q(bloque_in_1_57_) );
	DFFPOSX1 DFFPOSX1_727 ( .CLK(clk_bF_buf71), .D(_257__58_), .Q(bloque_in_1_58_) );
	DFFPOSX1 DFFPOSX1_728 ( .CLK(clk_bF_buf70), .D(_257__59_), .Q(bloque_in_1_59_) );
	DFFPOSX1 DFFPOSX1_729 ( .CLK(clk_bF_buf69), .D(_257__60_), .Q(bloque_in_1_60_) );
	DFFPOSX1 DFFPOSX1_730 ( .CLK(clk_bF_buf68), .D(_257__61_), .Q(bloque_in_1_61_) );
	DFFPOSX1 DFFPOSX1_731 ( .CLK(clk_bF_buf67), .D(_257__62_), .Q(bloque_in_1_62_) );
	DFFPOSX1 DFFPOSX1_732 ( .CLK(clk_bF_buf66), .D(_257__63_), .Q(bloque_in_1_63_) );
	DFFPOSX1 DFFPOSX1_733 ( .CLK(clk_bF_buf65), .D(_257__64_), .Q(bloque_in_1_64_) );
	DFFPOSX1 DFFPOSX1_734 ( .CLK(clk_bF_buf64), .D(_257__65_), .Q(bloque_in_1_65_) );
	DFFPOSX1 DFFPOSX1_735 ( .CLK(clk_bF_buf63), .D(_257__66_), .Q(bloque_in_1_66_) );
	DFFPOSX1 DFFPOSX1_736 ( .CLK(clk_bF_buf62), .D(_257__67_), .Q(bloque_in_1_67_) );
	DFFPOSX1 DFFPOSX1_737 ( .CLK(clk_bF_buf61), .D(_257__68_), .Q(bloque_in_1_68_) );
	DFFPOSX1 DFFPOSX1_738 ( .CLK(clk_bF_buf60), .D(_257__69_), .Q(bloque_in_1_69_) );
	DFFPOSX1 DFFPOSX1_739 ( .CLK(clk_bF_buf59), .D(_257__70_), .Q(bloque_in_1_70_) );
	DFFPOSX1 DFFPOSX1_740 ( .CLK(clk_bF_buf58), .D(_257__71_), .Q(bloque_in_1_71_) );
	DFFPOSX1 DFFPOSX1_741 ( .CLK(clk_bF_buf57), .D(_257__72_), .Q(bloque_in_1_72_) );
	DFFPOSX1 DFFPOSX1_742 ( .CLK(clk_bF_buf56), .D(_257__73_), .Q(bloque_in_1_73_) );
	DFFPOSX1 DFFPOSX1_743 ( .CLK(clk_bF_buf55), .D(_257__74_), .Q(bloque_in_1_74_) );
	DFFPOSX1 DFFPOSX1_744 ( .CLK(clk_bF_buf54), .D(_257__75_), .Q(bloque_in_1_75_) );
	DFFPOSX1 DFFPOSX1_745 ( .CLK(clk_bF_buf53), .D(_257__76_), .Q(bloque_in_1_76_) );
	DFFPOSX1 DFFPOSX1_746 ( .CLK(clk_bF_buf52), .D(_257__77_), .Q(bloque_in_1_77_) );
	DFFPOSX1 DFFPOSX1_747 ( .CLK(clk_bF_buf51), .D(_257__78_), .Q(bloque_in_1_78_) );
	DFFPOSX1 DFFPOSX1_748 ( .CLK(clk_bF_buf50), .D(_257__79_), .Q(bloque_in_1_79_) );
	DFFPOSX1 DFFPOSX1_749 ( .CLK(clk_bF_buf49), .D(_257__80_), .Q(bloque_in_1_80_) );
	DFFPOSX1 DFFPOSX1_750 ( .CLK(clk_bF_buf48), .D(_257__81_), .Q(bloque_in_1_81_) );
	DFFPOSX1 DFFPOSX1_751 ( .CLK(clk_bF_buf47), .D(_257__82_), .Q(bloque_in_1_82_) );
	DFFPOSX1 DFFPOSX1_752 ( .CLK(clk_bF_buf46), .D(_257__83_), .Q(bloque_in_1_83_) );
	DFFPOSX1 DFFPOSX1_753 ( .CLK(clk_bF_buf45), .D(_257__84_), .Q(bloque_in_1_84_) );
	DFFPOSX1 DFFPOSX1_754 ( .CLK(clk_bF_buf44), .D(_257__85_), .Q(bloque_in_1_85_) );
	DFFPOSX1 DFFPOSX1_755 ( .CLK(clk_bF_buf43), .D(_257__86_), .Q(bloque_in_1_86_) );
	DFFPOSX1 DFFPOSX1_756 ( .CLK(clk_bF_buf42), .D(_257__87_), .Q(bloque_in_1_87_) );
	DFFPOSX1 DFFPOSX1_757 ( .CLK(clk_bF_buf41), .D(_257__88_), .Q(bloque_in_1_88_) );
	DFFPOSX1 DFFPOSX1_758 ( .CLK(clk_bF_buf40), .D(_257__89_), .Q(bloque_in_1_89_) );
	DFFPOSX1 DFFPOSX1_759 ( .CLK(clk_bF_buf39), .D(_257__90_), .Q(bloque_in_1_90_) );
	DFFPOSX1 DFFPOSX1_760 ( .CLK(clk_bF_buf38), .D(_257__91_), .Q(bloque_in_1_91_) );
	DFFPOSX1 DFFPOSX1_761 ( .CLK(clk_bF_buf37), .D(_257__92_), .Q(bloque_in_1_92_) );
	DFFPOSX1 DFFPOSX1_762 ( .CLK(clk_bF_buf36), .D(_257__93_), .Q(bloque_in_1_93_) );
	DFFPOSX1 DFFPOSX1_763 ( .CLK(clk_bF_buf35), .D(_257__94_), .Q(bloque_in_1_94_) );
	DFFPOSX1 DFFPOSX1_764 ( .CLK(clk_bF_buf34), .D(_257__95_), .Q(bloque_in_1_95_) );
	DFFPOSX1 DFFPOSX1_765 ( .CLK(clk_bF_buf33), .D(_257__96_), .Q(bloque_in_1_96_) );
	DFFPOSX1 DFFPOSX1_766 ( .CLK(clk_bF_buf32), .D(_257__97_), .Q(bloque_in_1_97_) );
	DFFPOSX1 DFFPOSX1_767 ( .CLK(clk_bF_buf31), .D(_257__98_), .Q(bloque_in_1_98_) );
	DFFPOSX1 DFFPOSX1_768 ( .CLK(clk_bF_buf30), .D(_257__99_), .Q(bloque_in_1_99_) );
	DFFPOSX1 DFFPOSX1_769 ( .CLK(clk_bF_buf29), .D(_257__100_), .Q(bloque_in_1_100_) );
	DFFPOSX1 DFFPOSX1_770 ( .CLK(clk_bF_buf28), .D(_257__101_), .Q(bloque_in_1_101_) );
	DFFPOSX1 DFFPOSX1_771 ( .CLK(clk_bF_buf27), .D(_257__102_), .Q(bloque_in_1_102_) );
	DFFPOSX1 DFFPOSX1_772 ( .CLK(clk_bF_buf26), .D(_257__103_), .Q(bloque_in_1_103_) );
	DFFPOSX1 DFFPOSX1_773 ( .CLK(clk_bF_buf25), .D(_257__104_), .Q(bloque_in_1_104_) );
	DFFPOSX1 DFFPOSX1_774 ( .CLK(clk_bF_buf24), .D(_257__105_), .Q(bloque_in_1_105_) );
	DFFPOSX1 DFFPOSX1_775 ( .CLK(clk_bF_buf23), .D(_257__106_), .Q(bloque_in_1_106_) );
	DFFPOSX1 DFFPOSX1_776 ( .CLK(clk_bF_buf22), .D(_257__107_), .Q(bloque_in_1_107_) );
	DFFPOSX1 DFFPOSX1_777 ( .CLK(clk_bF_buf21), .D(_257__108_), .Q(bloque_in_1_108_) );
	DFFPOSX1 DFFPOSX1_778 ( .CLK(clk_bF_buf20), .D(_257__109_), .Q(bloque_in_1_109_) );
	DFFPOSX1 DFFPOSX1_779 ( .CLK(clk_bF_buf19), .D(_257__110_), .Q(bloque_in_1_110_) );
	DFFPOSX1 DFFPOSX1_780 ( .CLK(clk_bF_buf18), .D(_257__111_), .Q(bloque_in_1_111_) );
	DFFPOSX1 DFFPOSX1_781 ( .CLK(clk_bF_buf17), .D(_257__112_), .Q(bloque_in_1_112_) );
	DFFPOSX1 DFFPOSX1_782 ( .CLK(clk_bF_buf16), .D(_257__113_), .Q(bloque_in_1_113_) );
	DFFPOSX1 DFFPOSX1_783 ( .CLK(clk_bF_buf15), .D(_257__114_), .Q(bloque_in_1_114_) );
	DFFPOSX1 DFFPOSX1_784 ( .CLK(clk_bF_buf14), .D(_257__115_), .Q(bloque_in_1_115_) );
	DFFPOSX1 DFFPOSX1_785 ( .CLK(clk_bF_buf13), .D(_257__116_), .Q(bloque_in_1_116_) );
	DFFPOSX1 DFFPOSX1_786 ( .CLK(clk_bF_buf12), .D(_257__117_), .Q(bloque_in_1_117_) );
	DFFPOSX1 DFFPOSX1_787 ( .CLK(clk_bF_buf11), .D(_257__118_), .Q(bloque_in_1_118_) );
	DFFPOSX1 DFFPOSX1_788 ( .CLK(clk_bF_buf10), .D(_257__119_), .Q(bloque_in_1_119_) );
	DFFPOSX1 DFFPOSX1_789 ( .CLK(clk_bF_buf9), .D(_257__120_), .Q(bloque_in_1_120_) );
	DFFPOSX1 DFFPOSX1_790 ( .CLK(clk_bF_buf8), .D(_257__121_), .Q(bloque_in_1_121_) );
	DFFPOSX1 DFFPOSX1_791 ( .CLK(clk_bF_buf7), .D(_257__122_), .Q(bloque_in_1_122_) );
	DFFPOSX1 DFFPOSX1_792 ( .CLK(clk_bF_buf6), .D(_257__123_), .Q(bloque_in_1_123_) );
	DFFPOSX1 DFFPOSX1_793 ( .CLK(clk_bF_buf5), .D(_257__124_), .Q(bloque_in_1_124_) );
	DFFPOSX1 DFFPOSX1_794 ( .CLK(clk_bF_buf4), .D(_257__125_), .Q(bloque_in_1_125_) );
	DFFPOSX1 DFFPOSX1_795 ( .CLK(clk_bF_buf3), .D(_257__126_), .Q(bloque_in_1_126_) );
	DFFPOSX1 DFFPOSX1_796 ( .CLK(clk_bF_buf2), .D(_257__127_), .Q(bloque_in_1_127_) );
	INVX2 INVX2_3 ( .A(concatenador_counter_5_), .Y(_779_) );
	NOR2X1 NOR2X1_215 ( .A(concatenador_counter_1_bF_buf4), .B(_779_), .Y(_780_) );
	NOR3X1 NOR3X1_4 ( .A(concatenador_counter_4_), .B(concatenador_counter_3_), .C(concatenador_counter_2_), .Y(_781_) );
	NAND3X1 NAND3X1_123 ( .A(concatenador_counter_0_bF_buf10), .B(_781_), .C(_780_), .Y(_782_) );
	NAND2X1 NAND2X1_341 ( .A(reset_L_bF_buf36), .B(_782_), .Y(_783_) );
	OR2X2 OR2X2_21 ( .A(concatenador_counter_3_), .B(concatenador_counter_2_), .Y(_784_) );
	INVX1 INVX1_579 ( .A(concatenador_counter_1_bF_buf3), .Y(_785_) );
	INVX1 INVX1_580 ( .A(concatenador_counter_4_), .Y(_786_) );
	NAND3X1 NAND3X1_124 ( .A(concatenador_counter_5_), .B(_785_), .C(_786_), .Y(_787_) );
	NOR2X1 NOR2X1_216 ( .A(_784_), .B(_787_), .Y(_788_) );
	OAI21X1 OAI21X1_722 ( .A(_788_), .B(concatenador_counter_5_), .C(concatenador_counter_0_bF_buf9), .Y(_789_) );
	INVX1 INVX1_581 ( .A(concatenador_counter_0_bF_buf8), .Y(_790_) );
	OAI21X1 OAI21X1_723 ( .A(_788_), .B(_779_), .C(_790_), .Y(_791_) );
	AOI21X1 AOI21X1_575 ( .A(_789_), .B(_791_), .C(_783_), .Y(_778__0_) );
	AOI21X1 AOI21X1_576 ( .A(concatenador_counter_0_bF_buf7), .B(_779_), .C(concatenador_counter_1_bF_buf2), .Y(_792_) );
	NAND3X1 NAND3X1_125 ( .A(concatenador_counter_1_bF_buf1), .B(concatenador_counter_0_bF_buf6), .C(_779_), .Y(_793_) );
	NAND3X1 NAND3X1_126 ( .A(reset_L_bF_buf35), .B(_793_), .C(_782_), .Y(_794_) );
	NOR2X1 NOR2X1_217 ( .A(_792_), .B(_794_), .Y(_778__1_) );
	OAI21X1 OAI21X1_724 ( .A(_787_), .B(_784_), .C(concatenador_counter_5_), .Y(_795_) );
	NAND2X1 NAND2X1_342 ( .A(concatenador_counter_1_bF_buf0), .B(concatenador_counter_0_bF_buf5), .Y(_796_) );
	XNOR2X1 XNOR2X1_13 ( .A(_796_), .B(concatenador_counter_2_), .Y(_797_) );
	NAND3X1 NAND3X1_127 ( .A(_782_), .B(_797_), .C(_795_), .Y(_798_) );
	NAND2X1 NAND2X1_343 ( .A(concatenador_counter_5_), .B(_786_), .Y(_799_) );
	NAND2X1 NAND2X1_344 ( .A(concatenador_counter_0_bF_buf4), .B(_785_), .Y(_800_) );
	NOR3X1 NOR3X1_5 ( .A(_799_), .B(_784_), .C(_800_), .Y(_801_) );
	AOI21X1 AOI21X1_577 ( .A(_785_), .B(_781_), .C(_779_), .Y(_802_) );
	OAI21X1 OAI21X1_725 ( .A(_801_), .B(_802_), .C(concatenador_counter_2_), .Y(_803_) );
	AOI21X1 AOI21X1_578 ( .A(_798_), .B(_803_), .C(_783_), .Y(_778__2_) );
	NAND3X1 NAND3X1_128 ( .A(concatenador_counter_1_bF_buf7), .B(concatenador_counter_0_bF_buf3), .C(concatenador_counter_2_), .Y(_804_) );
	XNOR2X1 XNOR2X1_14 ( .A(_804_), .B(concatenador_counter_3_), .Y(_805_) );
	NAND3X1 NAND3X1_129 ( .A(_782_), .B(_805_), .C(_795_), .Y(_806_) );
	OAI21X1 OAI21X1_726 ( .A(_801_), .B(_802_), .C(concatenador_counter_3_), .Y(_807_) );
	AOI21X1 AOI21X1_579 ( .A(_806_), .B(_807_), .C(_783_), .Y(_778__3_) );
	NAND2X1 NAND2X1_345 ( .A(concatenador_counter_3_), .B(concatenador_counter_2_), .Y(_808_) );
	NOR2X1 NOR2X1_218 ( .A(_796_), .B(_808_), .Y(_809_) );
	NAND3X1 NAND3X1_130 ( .A(_782_), .B(_809_), .C(_795_), .Y(_810_) );
	NAND3X1 NAND3X1_131 ( .A(_779_), .B(concatenador_counter_4_), .C(_809_), .Y(_811_) );
	NAND3X1 NAND3X1_132 ( .A(reset_L_bF_buf34), .B(_782_), .C(_811_), .Y(_812_) );
	AOI21X1 AOI21X1_580 ( .A(_786_), .B(_810_), .C(_812_), .Y(_778__4_) );
	AOI21X1 AOI21X1_581 ( .A(_779_), .B(_811_), .C(_783_), .Y(_778__5_) );
	DFFPOSX1 DFFPOSX1_797 ( .CLK(clk_bF_buf1), .D(_778__0_), .Q(concatenador_counter_0_) );
	DFFPOSX1 DFFPOSX1_798 ( .CLK(clk_bF_buf0), .D(_778__1_), .Q(concatenador_counter_1_) );
	DFFPOSX1 DFFPOSX1_799 ( .CLK(clk_bF_buf113), .D(_778__2_), .Q(concatenador_counter_2_) );
	DFFPOSX1 DFFPOSX1_800 ( .CLK(clk_bF_buf112), .D(_778__3_), .Q(concatenador_counter_3_) );
	DFFPOSX1 DFFPOSX1_801 ( .CLK(clk_bF_buf111), .D(_778__4_), .Q(concatenador_counter_4_) );
	DFFPOSX1 DFFPOSX1_802 ( .CLK(clk_bF_buf110), .D(_778__5_), .Q(concatenador_counter_5_) );
	INVX1 INVX1_582 ( .A(concatenador_counter_0_bF_buf2), .Y(_815_) );
	NAND2X1 NAND2X1_346 ( .A(reset_L_bF_buf33), .B(_815_), .Y(_814__0_) );
	INVX1 INVX1_583 ( .A(concatenador_counter_1_bF_buf6), .Y(_816_) );
	NAND2X1 NAND2X1_347 ( .A(reset_L_bF_buf32), .B(_816_), .Y(_814__1_) );
	INVX1 INVX1_584 ( .A(concatenador_counter_2_), .Y(_817_) );
	NAND2X1 NAND2X1_348 ( .A(reset_L_bF_buf31), .B(_817_), .Y(_814__2_) );
	INVX1 INVX1_585 ( .A(concatenador_counter_3_), .Y(_818_) );
	NAND2X1 NAND2X1_349 ( .A(reset_L_bF_buf30), .B(_818_), .Y(_814__3_) );
	INVX1 INVX1_586 ( .A(concatenador_counter_4_), .Y(_819_) );
	NAND2X1 NAND2X1_350 ( .A(reset_L_bF_buf29), .B(_819_), .Y(_814__4_) );
	INVX1 INVX1_587 ( .A(concatenador_counter_5_), .Y(_820_) );
	NAND2X1 NAND2X1_351 ( .A(reset_L_bF_buf28), .B(_820_), .Y(_814__5_) );
	INVX1 INVX1_588 ( .A(contador_hash_synth_2_counter_d_0_), .Y(_821_) );
	NAND2X1 NAND2X1_352 ( .A(reset_L_bF_buf27), .B(_821_), .Y(_813__0_) );
	INVX1 INVX1_589 ( .A(contador_hash_synth_2_counter_d_1_), .Y(_822_) );
	NAND2X1 NAND2X1_353 ( .A(reset_L_bF_buf26), .B(_822_), .Y(_813__1_) );
	INVX1 INVX1_590 ( .A(contador_hash_synth_2_counter_d_2_), .Y(_823_) );
	NAND2X1 NAND2X1_354 ( .A(reset_L_bF_buf25), .B(_823_), .Y(_813__2_) );
	INVX1 INVX1_591 ( .A(contador_hash_synth_2_counter_d_3_), .Y(_824_) );
	NAND2X1 NAND2X1_355 ( .A(reset_L_bF_buf24), .B(_824_), .Y(_813__3_) );
	INVX1 INVX1_592 ( .A(contador_hash_synth_2_counter_d_4_), .Y(_825_) );
	NAND2X1 NAND2X1_356 ( .A(reset_L_bF_buf23), .B(_825_), .Y(_813__4_) );
	INVX1 INVX1_593 ( .A(contador_hash_synth_2_counter_d_5_), .Y(_826_) );
	NAND2X1 NAND2X1_357 ( .A(reset_L_bF_buf22), .B(_826_), .Y(_813__5_) );
	DFFPOSX1 DFFPOSX1_803 ( .CLK(clk_bF_buf109), .D(_813__0_), .Q(concatenador_counter_2d_0_) );
	DFFPOSX1 DFFPOSX1_804 ( .CLK(clk_bF_buf108), .D(_813__1_), .Q(concatenador_counter_2d_1_) );
	DFFPOSX1 DFFPOSX1_805 ( .CLK(clk_bF_buf107), .D(_813__2_), .Q(concatenador_counter_2d_2_) );
	DFFPOSX1 DFFPOSX1_806 ( .CLK(clk_bF_buf106), .D(_813__3_), .Q(concatenador_counter_2d_3_) );
	DFFPOSX1 DFFPOSX1_807 ( .CLK(clk_bF_buf105), .D(_813__4_), .Q(concatenador_counter_2d_4_) );
	DFFPOSX1 DFFPOSX1_808 ( .CLK(clk_bF_buf104), .D(_813__5_), .Q(concatenador_counter_2d_5_) );
	DFFPOSX1 DFFPOSX1_809 ( .CLK(clk_bF_buf103), .D(_814__0_), .Q(contador_hash_synth_2_counter_d_0_) );
	DFFPOSX1 DFFPOSX1_810 ( .CLK(clk_bF_buf102), .D(_814__1_), .Q(contador_hash_synth_2_counter_d_1_) );
	DFFPOSX1 DFFPOSX1_811 ( .CLK(clk_bF_buf101), .D(_814__2_), .Q(contador_hash_synth_2_counter_d_2_) );
	DFFPOSX1 DFFPOSX1_812 ( .CLK(clk_bF_buf100), .D(_814__3_), .Q(contador_hash_synth_2_counter_d_3_) );
	DFFPOSX1 DFFPOSX1_813 ( .CLK(clk_bF_buf99), .D(_814__4_), .Q(contador_hash_synth_2_counter_d_4_) );
	DFFPOSX1 DFFPOSX1_814 ( .CLK(clk_bF_buf98), .D(_814__5_), .Q(contador_hash_synth_2_counter_d_5_) );
	NOR2X1 NOR2X1_219 ( .A(reset_L_bF_buf21), .B(_1__bF_buf4), .Y(_829_) );
	INVX2 INVX2_4 ( .A(_829_), .Y(_830_) );
	AND2X2 AND2X2_33 ( .A(_830_), .B(gen_nonce_synth_rand_0_), .Y(_828__0_) );
	OR2X2 OR2X2_22 ( .A(_829_), .B(gen_nonce_synth_rand_1_), .Y(_828__1_) );
	INVX1 INVX1_594 ( .A(gen_nonce_synth_rand_2_), .Y(_831_) );
	NOR2X1 NOR2X1_220 ( .A(_831_), .B(_829_), .Y(_828__2_) );
	INVX1 INVX1_595 ( .A(gen_nonce_synth_rand_3_), .Y(_832_) );
	OAI21X1 OAI21X1_727 ( .A(reset_L_bF_buf20), .B(_1__bF_buf3), .C(_832_), .Y(_828__3_) );
	AND2X2 AND2X2_34 ( .A(_830_), .B(gen_nonce_synth_rand_4_), .Y(_828__4_) );
	AND2X2 AND2X2_35 ( .A(_830_), .B(gen_nonce_synth_rand_5_), .Y(_828__5_) );
	INVX1 INVX1_596 ( .A(gen_nonce_synth_rand_6_), .Y(_833_) );
	OAI21X1 OAI21X1_728 ( .A(reset_L_bF_buf19), .B(_1__bF_buf2), .C(_833_), .Y(_828__6_) );
	AND2X2 AND2X2_36 ( .A(_830_), .B(gen_nonce_synth_rand_7_), .Y(_828__7_) );
	INVX1 INVX1_597 ( .A(gen_nonce_synth_rand_8_), .Y(_834_) );
	NOR2X1 NOR2X1_221 ( .A(_834_), .B(_829_), .Y(_828__8_) );
	INVX1 INVX1_598 ( .A(gen_nonce_synth_rand_9_), .Y(_835_) );
	OAI21X1 OAI21X1_729 ( .A(reset_L_bF_buf18), .B(_1__bF_buf1), .C(_835_), .Y(_828__9_) );
	INVX1 INVX1_599 ( .A(gen_nonce_synth_rand_10_), .Y(_836_) );
	NOR2X1 NOR2X1_222 ( .A(_836_), .B(_829_), .Y(_828__10_) );
	INVX1 INVX1_600 ( .A(gen_nonce_synth_rand_11_), .Y(_837_) );
	NOR2X1 NOR2X1_223 ( .A(_837_), .B(_829_), .Y(_828__11_) );
	INVX1 INVX1_601 ( .A(gen_nonce_synth_rand_12_), .Y(_838_) );
	OAI21X1 OAI21X1_730 ( .A(reset_L_bF_buf17), .B(_1__bF_buf0), .C(_838_), .Y(_828__12_) );
	INVX1 INVX1_602 ( .A(gen_nonce_synth_rand_13_), .Y(_839_) );
	OAI21X1 OAI21X1_731 ( .A(reset_L_bF_buf16), .B(_1__bF_buf5), .C(_839_), .Y(_828__13_) );
	INVX1 INVX1_603 ( .A(gen_nonce_synth_rand_14_), .Y(_840_) );
	OAI21X1 OAI21X1_732 ( .A(reset_L_bF_buf15), .B(_1__bF_buf4), .C(_840_), .Y(_828__14_) );
	INVX1 INVX1_604 ( .A(gen_nonce_synth_rand_15_), .Y(_841_) );
	NOR2X1 NOR2X1_224 ( .A(_841_), .B(_829_), .Y(_828__15_) );
	INVX1 INVX1_605 ( .A(gen_nonce_synth_rand_16_), .Y(_842_) );
	OAI21X1 OAI21X1_733 ( .A(reset_L_bF_buf14), .B(_1__bF_buf3), .C(_842_), .Y(_828__16_) );
	INVX1 INVX1_606 ( .A(gen_nonce_synth_rand_17_), .Y(_843_) );
	OAI21X1 OAI21X1_734 ( .A(reset_L_bF_buf13), .B(_1__bF_buf2), .C(_843_), .Y(_828__17_) );
	INVX1 INVX1_607 ( .A(gen_nonce_synth_rand_18_), .Y(_844_) );
	NOR2X1 NOR2X1_225 ( .A(_844_), .B(_829_), .Y(_828__18_) );
	INVX1 INVX1_608 ( .A(gen_nonce_synth_rand_19_), .Y(_845_) );
	OAI21X1 OAI21X1_735 ( .A(reset_L_bF_buf12), .B(_1__bF_buf1), .C(_845_), .Y(_828__19_) );
	INVX1 INVX1_609 ( .A(gen_nonce_synth_rand_20_), .Y(_846_) );
	NOR2X1 NOR2X1_226 ( .A(_846_), .B(_829_), .Y(_828__20_) );
	INVX1 INVX1_610 ( .A(gen_nonce_synth_rand_21_), .Y(_847_) );
	NOR2X1 NOR2X1_227 ( .A(_847_), .B(_829_), .Y(_828__21_) );
	INVX1 INVX1_611 ( .A(gen_nonce_synth_rand_22_), .Y(_848_) );
	OAI21X1 OAI21X1_736 ( .A(reset_L_bF_buf11), .B(_1__bF_buf0), .C(_848_), .Y(_828__22_) );
	INVX1 INVX1_612 ( .A(gen_nonce_synth_rand_23_), .Y(_849_) );
	NOR2X1 NOR2X1_228 ( .A(_849_), .B(_829_), .Y(_828__23_) );
	INVX1 INVX1_613 ( .A(gen_nonce_synth_rand_24_), .Y(_850_) );
	OAI21X1 OAI21X1_737 ( .A(reset_L_bF_buf10), .B(_1__bF_buf5), .C(_850_), .Y(_828__24_) );
	INVX1 INVX1_614 ( .A(gen_nonce_synth_rand_25_), .Y(_851_) );
	OAI21X1 OAI21X1_738 ( .A(reset_L_bF_buf9), .B(_1__bF_buf4), .C(_851_), .Y(_828__25_) );
	AND2X2 AND2X2_37 ( .A(_830_), .B(gen_nonce_synth_rand_26_), .Y(_828__26_) );
	AND2X2 AND2X2_38 ( .A(_830_), .B(gen_nonce_synth_rand_27_), .Y(_828__27_) );
	INVX1 INVX1_615 ( .A(gen_nonce_synth_rand_28_), .Y(_852_) );
	NOR2X1 NOR2X1_229 ( .A(_852_), .B(_829_), .Y(_828__28_) );
	INVX1 INVX1_616 ( .A(gen_nonce_synth_rand_29_), .Y(_853_) );
	OAI21X1 OAI21X1_739 ( .A(reset_L_bF_buf8), .B(_1__bF_buf3), .C(_853_), .Y(_828__29_) );
	AND2X2 AND2X2_39 ( .A(_830_), .B(gen_nonce_synth_rand_30_), .Y(_828__30_) );
	AND2X2 AND2X2_40 ( .A(_830_), .B(gen_nonce_synth_rand_31_), .Y(_828__31_) );
	INVX4 INVX4_2 ( .A(_1__bF_buf2), .Y(_854_) );
	INVX8 INVX8_5 ( .A(comparador_valid_bF_buf1), .Y(_855_) );
	NAND3X1 NAND3X1_133 ( .A(gen_nonce_synth_rand_0_), .B(_854_), .C(_855__bF_buf4), .Y(_856_) );
	AND2X2 AND2X2_41 ( .A(_856_), .B(_2__0_), .Y(_857_) );
	OAI21X1 OAI21X1_740 ( .A(_856_), .B(_2__0_), .C(_830_), .Y(_858_) );
	OR2X2 OR2X2_23 ( .A(_857_), .B(_858_), .Y(_827__0_) );
	INVX1 INVX1_617 ( .A(_2__1_), .Y(_859_) );
	NAND2X1 NAND2X1_358 ( .A(gen_nonce_synth_rand_0_), .B(_2__0_), .Y(_860_) );
	AND2X2 AND2X2_42 ( .A(gen_nonce_synth_rand_1_), .B(_2__1_), .Y(_861_) );
	NOR2X1 NOR2X1_230 ( .A(gen_nonce_synth_rand_1_), .B(_2__1_), .Y(_862_) );
	NOR2X1 NOR2X1_231 ( .A(_862_), .B(_861_), .Y(_863_) );
	XNOR2X1 XNOR2X1_15 ( .A(_863_), .B(_860_), .Y(_864_) );
	NAND2X1 NAND2X1_359 ( .A(comparador_valid_bF_buf0), .B(_859_), .Y(_865_) );
	OAI21X1 OAI21X1_741 ( .A(_864_), .B(comparador_valid_bF_buf5), .C(_865_), .Y(_866_) );
	NAND2X1 NAND2X1_360 ( .A(reset_L_bF_buf7), .B(_854_), .Y(_867_) );
	INVX4 INVX4_3 ( .A(_867_), .Y(_868_) );
	AOI22X1 AOI22X1_14 ( .A(_1__bF_buf1), .B(_859_), .C(_866_), .D(_868__bF_buf3), .Y(_827__1_) );
	INVX1 INVX1_618 ( .A(_2__2_), .Y(_869_) );
	AND2X2 AND2X2_43 ( .A(gen_nonce_synth_rand_0_), .B(_2__0_), .Y(_870_) );
	OR2X2 OR2X2_24 ( .A(gen_nonce_synth_rand_1_), .B(_2__1_), .Y(_871_) );
	AOI21X1 AOI21X1_582 ( .A(_870_), .B(_871_), .C(_861_), .Y(_872_) );
	XNOR2X1 XNOR2X1_16 ( .A(gen_nonce_synth_rand_2_), .B(_2__2_), .Y(_873_) );
	NOR2X1 NOR2X1_232 ( .A(_873_), .B(_872_), .Y(_874_) );
	AND2X2 AND2X2_44 ( .A(_872_), .B(_873_), .Y(_875_) );
	OAI21X1 OAI21X1_742 ( .A(_875_), .B(_874_), .C(_855__bF_buf3), .Y(_876_) );
	OAI21X1 OAI21X1_743 ( .A(_855__bF_buf2), .B(_2__2_), .C(_876_), .Y(_877_) );
	AOI22X1 AOI22X1_15 ( .A(_1__bF_buf0), .B(_869_), .C(_877_), .D(_868__bF_buf2), .Y(_827__2_) );
	INVX1 INVX1_619 ( .A(_2__3_), .Y(_878_) );
	XNOR2X1 XNOR2X1_17 ( .A(gen_nonce_synth_rand_3_), .B(_2__3_), .Y(_879_) );
	NAND2X1 NAND2X1_361 ( .A(gen_nonce_synth_rand_2_), .B(_2__2_), .Y(_880_) );
	OAI21X1 OAI21X1_744 ( .A(_872_), .B(_873_), .C(_880_), .Y(_881_) );
	OAI21X1 OAI21X1_745 ( .A(_881_), .B(_879_), .C(_855__bF_buf1), .Y(_882_) );
	AOI21X1 AOI21X1_583 ( .A(_879_), .B(_881_), .C(_882_), .Y(_883_) );
	OAI21X1 OAI21X1_746 ( .A(_855__bF_buf0), .B(_2__3_), .C(_868__bF_buf1), .Y(_884_) );
	OAI22X1 OAI22X1_219 ( .A(_854_), .B(_878_), .C(_883_), .D(_884_), .Y(_827__3_) );
	NAND2X1 NAND2X1_362 ( .A(_1__bF_buf5), .B(_2__4_), .Y(_885_) );
	INVX1 INVX1_620 ( .A(_861_), .Y(_886_) );
	OAI21X1 OAI21X1_747 ( .A(_862_), .B(_860_), .C(_886_), .Y(_887_) );
	NAND2X1 NAND2X1_363 ( .A(gen_nonce_synth_rand_2_), .B(_869_), .Y(_888_) );
	NAND2X1 NAND2X1_364 ( .A(_2__2_), .B(_831_), .Y(_889_) );
	NAND2X1 NAND2X1_365 ( .A(gen_nonce_synth_rand_3_), .B(_878_), .Y(_890_) );
	NAND2X1 NAND2X1_366 ( .A(_2__3_), .B(_832_), .Y(_891_) );
	AOI22X1 AOI22X1_16 ( .A(_888_), .B(_889_), .C(_890_), .D(_891_), .Y(_892_) );
	NAND2X1 NAND2X1_367 ( .A(gen_nonce_synth_rand_3_), .B(_2__3_), .Y(_893_) );
	NOR2X1 NOR2X1_233 ( .A(gen_nonce_synth_rand_3_), .B(_2__3_), .Y(_894_) );
	OAI21X1 OAI21X1_748 ( .A(_894_), .B(_880_), .C(_893_), .Y(_895_) );
	AOI21X1 AOI21X1_584 ( .A(_887_), .B(_892_), .C(_895_), .Y(_896_) );
	XNOR2X1 XNOR2X1_18 ( .A(gen_nonce_synth_rand_4_), .B(_2__4_), .Y(_897_) );
	NAND2X1 NAND2X1_368 ( .A(_897_), .B(_896_), .Y(_898_) );
	NOR3X1 NOR3X1_6 ( .A(_873_), .B(_879_), .C(_872_), .Y(_899_) );
	XOR2X1 XOR2X1_17 ( .A(gen_nonce_synth_rand_4_), .B(_2__4_), .Y(_900_) );
	OAI21X1 OAI21X1_749 ( .A(_899_), .B(_895_), .C(_900_), .Y(_901_) );
	AOI21X1 AOI21X1_585 ( .A(_898_), .B(_901_), .C(comparador_valid_bF_buf4), .Y(_902_) );
	OAI21X1 OAI21X1_750 ( .A(_855__bF_buf4), .B(_2__4_), .C(_868__bF_buf0), .Y(_903_) );
	OAI21X1 OAI21X1_751 ( .A(_902_), .B(_903_), .C(_885_), .Y(_827__4_) );
	NAND2X1 NAND2X1_369 ( .A(gen_nonce_synth_rand_4_), .B(_2__4_), .Y(_904_) );
	OAI21X1 OAI21X1_752 ( .A(_896_), .B(_897_), .C(_904_), .Y(_905_) );
	INVX1 INVX1_621 ( .A(_905_), .Y(_906_) );
	XNOR2X1 XNOR2X1_19 ( .A(gen_nonce_synth_rand_5_), .B(_2__5_), .Y(_907_) );
	AOI21X1 AOI21X1_586 ( .A(_907_), .B(_906_), .C(comparador_valid_bF_buf3), .Y(_908_) );
	OAI21X1 OAI21X1_753 ( .A(_906_), .B(_907_), .C(_908_), .Y(_909_) );
	AOI21X1 AOI21X1_587 ( .A(comparador_valid_bF_buf2), .B(_2__5_), .C(_867_), .Y(_910_) );
	NOR2X1 NOR2X1_234 ( .A(_2__5_), .B(_854_), .Y(_911_) );
	AOI21X1 AOI21X1_588 ( .A(_910_), .B(_909_), .C(_911_), .Y(_827__5_) );
	INVX1 INVX1_622 ( .A(_2__6_), .Y(_912_) );
	NAND2X1 NAND2X1_370 ( .A(gen_nonce_synth_rand_5_), .B(_2__5_), .Y(_913_) );
	NOR2X1 NOR2X1_235 ( .A(gen_nonce_synth_rand_5_), .B(_2__5_), .Y(_914_) );
	OAI21X1 OAI21X1_754 ( .A(_914_), .B(_904_), .C(_913_), .Y(_915_) );
	INVX1 INVX1_623 ( .A(_915_), .Y(_916_) );
	XOR2X1 XOR2X1_18 ( .A(gen_nonce_synth_rand_5_), .B(_2__5_), .Y(_917_) );
	NAND2X1 NAND2X1_371 ( .A(_900_), .B(_917_), .Y(_918_) );
	OAI21X1 OAI21X1_755 ( .A(_896_), .B(_918_), .C(_916_), .Y(_919_) );
	INVX1 INVX1_624 ( .A(_919_), .Y(_920_) );
	XNOR2X1 XNOR2X1_20 ( .A(gen_nonce_synth_rand_6_), .B(_2__6_), .Y(_921_) );
	AOI21X1 AOI21X1_589 ( .A(_921_), .B(_920_), .C(comparador_valid_bF_buf1), .Y(_922_) );
	OAI21X1 OAI21X1_756 ( .A(_920_), .B(_921_), .C(_922_), .Y(_923_) );
	AOI21X1 AOI21X1_590 ( .A(comparador_valid_bF_buf0), .B(_2__6_), .C(_867_), .Y(_924_) );
	AOI22X1 AOI22X1_17 ( .A(_1__bF_buf4), .B(_912_), .C(_923_), .D(_924_), .Y(_827__6_) );
	NAND2X1 NAND2X1_372 ( .A(gen_nonce_synth_rand_6_), .B(_2__6_), .Y(_925_) );
	OAI21X1 OAI21X1_757 ( .A(_920_), .B(_921_), .C(_925_), .Y(_926_) );
	XOR2X1 XOR2X1_19 ( .A(gen_nonce_synth_rand_7_), .B(_2__7_), .Y(_927_) );
	AND2X2 AND2X2_45 ( .A(_926_), .B(_927_), .Y(_928_) );
	OAI21X1 OAI21X1_758 ( .A(_926_), .B(_927_), .C(_855__bF_buf3), .Y(_929_) );
	AOI21X1 AOI21X1_591 ( .A(comparador_valid_bF_buf5), .B(_2__7_), .C(_867_), .Y(_930_) );
	OAI21X1 OAI21X1_759 ( .A(_928_), .B(_929_), .C(_930_), .Y(_931_) );
	OR2X2 OR2X2_25 ( .A(_854_), .B(_2__7_), .Y(_932_) );
	AND2X2 AND2X2_46 ( .A(_931_), .B(_932_), .Y(_827__7_) );
	INVX1 INVX1_625 ( .A(_2__8_), .Y(_933_) );
	NOR2X1 NOR2X1_236 ( .A(_897_), .B(_907_), .Y(_934_) );
	XNOR2X1 XNOR2X1_21 ( .A(gen_nonce_synth_rand_7_), .B(_2__7_), .Y(_935_) );
	NOR2X1 NOR2X1_237 ( .A(_921_), .B(_935_), .Y(_936_) );
	NAND2X1 NAND2X1_373 ( .A(_934_), .B(_936_), .Y(_937_) );
	NAND2X1 NAND2X1_374 ( .A(gen_nonce_synth_rand_7_), .B(_2__7_), .Y(_938_) );
	OAI21X1 OAI21X1_760 ( .A(_935_), .B(_925_), .C(_938_), .Y(_939_) );
	AOI21X1 AOI21X1_592 ( .A(_915_), .B(_936_), .C(_939_), .Y(_940_) );
	OAI21X1 OAI21X1_761 ( .A(_937_), .B(_896_), .C(_940_), .Y(_941_) );
	XOR2X1 XOR2X1_20 ( .A(gen_nonce_synth_rand_8_), .B(_2__8_), .Y(_942_) );
	NAND2X1 NAND2X1_375 ( .A(_942_), .B(_941_), .Y(_943_) );
	OR2X2 OR2X2_26 ( .A(_941_), .B(_942_), .Y(_944_) );
	NAND3X1 NAND3X1_134 ( .A(_855__bF_buf2), .B(_943_), .C(_944_), .Y(_945_) );
	AOI21X1 AOI21X1_593 ( .A(comparador_valid_bF_buf4), .B(_2__8_), .C(_867_), .Y(_946_) );
	AOI22X1 AOI22X1_18 ( .A(_1__bF_buf3), .B(_933_), .C(_945_), .D(_946_), .Y(_827__8_) );
	INVX1 INVX1_626 ( .A(_2__9_), .Y(_947_) );
	XOR2X1 XOR2X1_21 ( .A(gen_nonce_synth_rand_9_), .B(_2__9_), .Y(_948_) );
	INVX1 INVX1_627 ( .A(_948_), .Y(_949_) );
	OAI21X1 OAI21X1_762 ( .A(_834_), .B(_933_), .C(_943_), .Y(_950_) );
	OAI21X1 OAI21X1_763 ( .A(_950_), .B(_949_), .C(_855__bF_buf1), .Y(_951_) );
	AOI21X1 AOI21X1_594 ( .A(_949_), .B(_950_), .C(_951_), .Y(_952_) );
	OAI21X1 OAI21X1_764 ( .A(_855__bF_buf0), .B(_2__9_), .C(_868__bF_buf3), .Y(_953_) );
	OAI22X1 OAI22X1_220 ( .A(_854_), .B(_947_), .C(_952_), .D(_953_), .Y(_827__9_) );
	INVX1 INVX1_628 ( .A(_2__10_), .Y(_954_) );
	NOR2X1 NOR2X1_238 ( .A(_834_), .B(_933_), .Y(_955_) );
	NOR2X1 NOR2X1_239 ( .A(_835_), .B(_947_), .Y(_956_) );
	NAND2X1 NAND2X1_376 ( .A(_835_), .B(_947_), .Y(_957_) );
	OAI21X1 OAI21X1_765 ( .A(_955_), .B(_956_), .C(_957_), .Y(_958_) );
	OAI21X1 OAI21X1_766 ( .A(_943_), .B(_949_), .C(_958_), .Y(_959_) );
	XOR2X1 XOR2X1_22 ( .A(gen_nonce_synth_rand_10_), .B(_2__10_), .Y(_960_) );
	NAND2X1 NAND2X1_377 ( .A(_960_), .B(_959_), .Y(_961_) );
	INVX1 INVX1_629 ( .A(_959_), .Y(_962_) );
	INVX1 INVX1_630 ( .A(_960_), .Y(_963_) );
	NAND2X1 NAND2X1_378 ( .A(_963_), .B(_962_), .Y(_964_) );
	AOI21X1 AOI21X1_595 ( .A(_961_), .B(_964_), .C(comparador_valid_bF_buf3), .Y(_965_) );
	OAI21X1 OAI21X1_767 ( .A(_855__bF_buf4), .B(_2__10_), .C(_868__bF_buf2), .Y(_966_) );
	OAI22X1 OAI22X1_221 ( .A(_854_), .B(_954_), .C(_965_), .D(_966_), .Y(_827__10_) );
	INVX1 INVX1_631 ( .A(_2__11_), .Y(_967_) );
	OAI21X1 OAI21X1_768 ( .A(_836_), .B(_954_), .C(_961_), .Y(_968_) );
	XOR2X1 XOR2X1_23 ( .A(gen_nonce_synth_rand_11_), .B(_2__11_), .Y(_969_) );
	AND2X2 AND2X2_47 ( .A(_968_), .B(_969_), .Y(_970_) );
	OAI21X1 OAI21X1_769 ( .A(_968_), .B(_969_), .C(_855__bF_buf3), .Y(_971_) );
	OR2X2 OR2X2_27 ( .A(_970_), .B(_971_), .Y(_972_) );
	AOI21X1 AOI21X1_596 ( .A(comparador_valid_bF_buf2), .B(_2__11_), .C(_867_), .Y(_973_) );
	AOI22X1 AOI22X1_19 ( .A(_1__bF_buf2), .B(_967_), .C(_972_), .D(_973_), .Y(_827__11_) );
	NOR2X1 NOR2X1_240 ( .A(_2__12_), .B(_854_), .Y(_974_) );
	NOR2X1 NOR2X1_241 ( .A(_836_), .B(_954_), .Y(_975_) );
	NOR2X1 NOR2X1_242 ( .A(_837_), .B(_967_), .Y(_976_) );
	AOI21X1 AOI21X1_597 ( .A(_975_), .B(_969_), .C(_976_), .Y(_977_) );
	NAND2X1 NAND2X1_379 ( .A(_960_), .B(_969_), .Y(_978_) );
	OAI21X1 OAI21X1_770 ( .A(_978_), .B(_958_), .C(_977_), .Y(_979_) );
	NAND2X1 NAND2X1_380 ( .A(_942_), .B(_948_), .Y(_980_) );
	NOR2X1 NOR2X1_243 ( .A(_980_), .B(_978_), .Y(_981_) );
	AOI21X1 AOI21X1_598 ( .A(_981_), .B(_941_), .C(_979_), .Y(_982_) );
	XNOR2X1 XNOR2X1_22 ( .A(gen_nonce_synth_rand_12_), .B(_2__12_), .Y(_983_) );
	AOI21X1 AOI21X1_599 ( .A(_983_), .B(_982_), .C(comparador_valid_bF_buf1), .Y(_984_) );
	OAI21X1 OAI21X1_771 ( .A(_982_), .B(_983_), .C(_984_), .Y(_985_) );
	AOI21X1 AOI21X1_600 ( .A(comparador_valid_bF_buf0), .B(_2__12_), .C(_867_), .Y(_986_) );
	AOI21X1 AOI21X1_601 ( .A(_986_), .B(_985_), .C(_974_), .Y(_827__12_) );
	INVX1 INVX1_632 ( .A(_2__13_), .Y(_987_) );
	XNOR2X1 XNOR2X1_23 ( .A(gen_nonce_synth_rand_13_), .B(_2__13_), .Y(_988_) );
	NAND2X1 NAND2X1_381 ( .A(gen_nonce_synth_rand_12_), .B(_2__12_), .Y(_989_) );
	OAI21X1 OAI21X1_772 ( .A(_982_), .B(_983_), .C(_989_), .Y(_990_) );
	OAI21X1 OAI21X1_773 ( .A(_990_), .B(_988_), .C(_855__bF_buf2), .Y(_991_) );
	AOI21X1 AOI21X1_602 ( .A(_988_), .B(_990_), .C(_991_), .Y(_992_) );
	OAI21X1 OAI21X1_774 ( .A(_855__bF_buf1), .B(_2__13_), .C(_868__bF_buf1), .Y(_993_) );
	OAI22X1 OAI22X1_222 ( .A(_854_), .B(_987_), .C(_992_), .D(_993_), .Y(_827__13_) );
	INVX1 INVX1_633 ( .A(_2__14_), .Y(_994_) );
	XOR2X1 XOR2X1_24 ( .A(gen_nonce_synth_rand_12_), .B(_2__12_), .Y(_995_) );
	NAND2X1 NAND2X1_382 ( .A(gen_nonce_synth_rand_13_), .B(_2__13_), .Y(_996_) );
	NAND2X1 NAND2X1_383 ( .A(_839_), .B(_987_), .Y(_997_) );
	NAND3X1 NAND3X1_135 ( .A(_996_), .B(_997_), .C(_995_), .Y(_998_) );
	OAI21X1 OAI21X1_775 ( .A(_839_), .B(_987_), .C(_989_), .Y(_999_) );
	OAI21X1 OAI21X1_776 ( .A(gen_nonce_synth_rand_13_), .B(_2__13_), .C(_999_), .Y(_1000_) );
	OAI21X1 OAI21X1_777 ( .A(_982_), .B(_998_), .C(_1000_), .Y(_1001_) );
	XOR2X1 XOR2X1_25 ( .A(gen_nonce_synth_rand_14_), .B(_2__14_), .Y(_1002_) );
	AND2X2 AND2X2_48 ( .A(_1001_), .B(_1002_), .Y(_1003_) );
	OAI21X1 OAI21X1_778 ( .A(_1001_), .B(_1002_), .C(_855__bF_buf0), .Y(_1004_) );
	OR2X2 OR2X2_28 ( .A(_1003_), .B(_1004_), .Y(_1005_) );
	AOI21X1 AOI21X1_603 ( .A(comparador_valid_bF_buf5), .B(_2__14_), .C(_867_), .Y(_1006_) );
	AOI22X1 AOI22X1_20 ( .A(_1__bF_buf1), .B(_994_), .C(_1005_), .D(_1006_), .Y(_827__14_) );
	INVX1 INVX1_634 ( .A(_2__15_), .Y(_1007_) );
	NOR2X1 NOR2X1_244 ( .A(_840_), .B(_994_), .Y(_1008_) );
	NOR2X1 NOR2X1_245 ( .A(_1008_), .B(_1003_), .Y(_1009_) );
	XNOR2X1 XNOR2X1_24 ( .A(gen_nonce_synth_rand_15_), .B(_2__15_), .Y(_1010_) );
	AOI21X1 AOI21X1_604 ( .A(_1010_), .B(_1009_), .C(comparador_valid_bF_buf4), .Y(_1011_) );
	OAI21X1 OAI21X1_779 ( .A(_1009_), .B(_1010_), .C(_1011_), .Y(_1012_) );
	AOI21X1 AOI21X1_605 ( .A(comparador_valid_bF_buf3), .B(_2__15_), .C(_867_), .Y(_1013_) );
	AOI22X1 AOI22X1_21 ( .A(_1__bF_buf0), .B(_1007_), .C(_1012_), .D(_1013_), .Y(_827__15_) );
	INVX1 INVX1_635 ( .A(_2__16_), .Y(_1014_) );
	NOR2X1 NOR2X1_246 ( .A(_2__6_), .B(_833_), .Y(_1015_) );
	NOR2X1 NOR2X1_247 ( .A(gen_nonce_synth_rand_6_), .B(_912_), .Y(_1016_) );
	OAI21X1 OAI21X1_780 ( .A(_1015_), .B(_1016_), .C(_927_), .Y(_1017_) );
	NOR2X1 NOR2X1_248 ( .A(_918_), .B(_1017_), .Y(_1018_) );
	OAI21X1 OAI21X1_781 ( .A(_899_), .B(_895_), .C(_1018_), .Y(_1019_) );
	XOR2X1 XOR2X1_26 ( .A(gen_nonce_synth_rand_15_), .B(_2__15_), .Y(_1020_) );
	NAND2X1 NAND2X1_384 ( .A(_1002_), .B(_1020_), .Y(_1021_) );
	NOR2X1 NOR2X1_249 ( .A(_1021_), .B(_998_), .Y(_1022_) );
	NAND2X1 NAND2X1_385 ( .A(_981_), .B(_1022_), .Y(_1023_) );
	AOI21X1 AOI21X1_606 ( .A(_940_), .B(_1019_), .C(_1023_), .Y(_1024_) );
	NOR2X1 NOR2X1_250 ( .A(_841_), .B(_1007_), .Y(_1025_) );
	AOI21X1 AOI21X1_607 ( .A(_1008_), .B(_1020_), .C(_1025_), .Y(_1026_) );
	OAI21X1 OAI21X1_782 ( .A(_1021_), .B(_1000_), .C(_1026_), .Y(_1027_) );
	AOI21X1 AOI21X1_608 ( .A(_1022_), .B(_979_), .C(_1027_), .Y(_1028_) );
	INVX1 INVX1_636 ( .A(_1028_), .Y(_1029_) );
	NOR2X1 NOR2X1_251 ( .A(_1029_), .B(_1024_), .Y(_1030_) );
	NAND2X1 NAND2X1_386 ( .A(gen_nonce_synth_rand_16_), .B(_2__16_), .Y(_1031_) );
	NAND2X1 NAND2X1_387 ( .A(_842_), .B(_1014_), .Y(_1032_) );
	NAND2X1 NAND2X1_388 ( .A(_1031_), .B(_1032_), .Y(_1033_) );
	AOI21X1 AOI21X1_609 ( .A(_1033_), .B(_1030_), .C(comparador_valid_bF_buf2), .Y(_1034_) );
	OAI21X1 OAI21X1_783 ( .A(_1030_), .B(_1033_), .C(_1034_), .Y(_1035_) );
	AOI21X1 AOI21X1_610 ( .A(comparador_valid_bF_buf1), .B(_2__16_), .C(_867_), .Y(_1036_) );
	AOI22X1 AOI22X1_22 ( .A(_1__bF_buf5), .B(_1014_), .C(_1035_), .D(_1036_), .Y(_827__16_) );
	INVX1 INVX1_637 ( .A(_2__17_), .Y(_1037_) );
	OAI21X1 OAI21X1_784 ( .A(_1030_), .B(_1033_), .C(_1031_), .Y(_1038_) );
	NOR2X1 NOR2X1_252 ( .A(_843_), .B(_1037_), .Y(_1039_) );
	NOR2X1 NOR2X1_253 ( .A(gen_nonce_synth_rand_17_), .B(_2__17_), .Y(_1040_) );
	OR2X2 OR2X2_29 ( .A(_1039_), .B(_1040_), .Y(_1041_) );
	OAI21X1 OAI21X1_785 ( .A(_1038_), .B(_1041_), .C(_855__bF_buf4), .Y(_1042_) );
	AOI21X1 AOI21X1_611 ( .A(_1038_), .B(_1041_), .C(_1042_), .Y(_1043_) );
	OAI21X1 OAI21X1_786 ( .A(_855__bF_buf3), .B(_2__17_), .C(_868__bF_buf0), .Y(_1044_) );
	OAI22X1 OAI22X1_223 ( .A(_854_), .B(_1037_), .C(_1043_), .D(_1044_), .Y(_827__17_) );
	INVX1 INVX1_638 ( .A(_2__18_), .Y(_1045_) );
	OAI21X1 OAI21X1_787 ( .A(_843_), .B(_1037_), .C(_1031_), .Y(_1046_) );
	OAI21X1 OAI21X1_788 ( .A(gen_nonce_synth_rand_17_), .B(_2__17_), .C(_1046_), .Y(_1047_) );
	NOR2X1 NOR2X1_254 ( .A(_1033_), .B(_1041_), .Y(_1048_) );
	INVX1 INVX1_639 ( .A(_1048_), .Y(_1049_) );
	OAI21X1 OAI21X1_789 ( .A(_1030_), .B(_1049_), .C(_1047_), .Y(_1050_) );
	NAND2X1 NAND2X1_389 ( .A(gen_nonce_synth_rand_18_), .B(_2__18_), .Y(_1051_) );
	NAND2X1 NAND2X1_390 ( .A(_844_), .B(_1045_), .Y(_1052_) );
	AND2X2 AND2X2_49 ( .A(_1052_), .B(_1051_), .Y(_1053_) );
	OR2X2 OR2X2_30 ( .A(_1050_), .B(_1053_), .Y(_1054_) );
	NAND2X1 NAND2X1_391 ( .A(_1053_), .B(_1050_), .Y(_1055_) );
	AOI21X1 AOI21X1_612 ( .A(_1055_), .B(_1054_), .C(comparador_valid_bF_buf0), .Y(_1056_) );
	OAI21X1 OAI21X1_790 ( .A(_855__bF_buf2), .B(_2__18_), .C(_868__bF_buf3), .Y(_1057_) );
	OAI22X1 OAI22X1_224 ( .A(_854_), .B(_1045_), .C(_1056_), .D(_1057_), .Y(_827__18_) );
	INVX1 INVX1_640 ( .A(_2__19_), .Y(_1058_) );
	AND2X2 AND2X2_50 ( .A(_1055_), .B(_1051_), .Y(_1059_) );
	NAND2X1 NAND2X1_392 ( .A(gen_nonce_synth_rand_19_), .B(_2__19_), .Y(_1060_) );
	NAND2X1 NAND2X1_393 ( .A(_845_), .B(_1058_), .Y(_1061_) );
	NAND2X1 NAND2X1_394 ( .A(_1060_), .B(_1061_), .Y(_1062_) );
	AOI21X1 AOI21X1_613 ( .A(_1062_), .B(_1059_), .C(comparador_valid_bF_buf5), .Y(_1063_) );
	OAI21X1 OAI21X1_791 ( .A(_1059_), .B(_1062_), .C(_1063_), .Y(_1064_) );
	AOI21X1 AOI21X1_614 ( .A(comparador_valid_bF_buf4), .B(_2__19_), .C(_867_), .Y(_1065_) );
	AOI22X1 AOI22X1_23 ( .A(_1__bF_buf4), .B(_1058_), .C(_1064_), .D(_1065_), .Y(_827__19_) );
	INVX1 INVX1_641 ( .A(_2__20_), .Y(_1066_) );
	INVX1 INVX1_642 ( .A(_1047_), .Y(_1067_) );
	NAND2X1 NAND2X1_395 ( .A(_1051_), .B(_1052_), .Y(_1068_) );
	NOR2X1 NOR2X1_255 ( .A(_1068_), .B(_1062_), .Y(_1069_) );
	OAI21X1 OAI21X1_792 ( .A(_1062_), .B(_1051_), .C(_1060_), .Y(_1070_) );
	AOI21X1 AOI21X1_615 ( .A(_1069_), .B(_1067_), .C(_1070_), .Y(_1071_) );
	NAND2X1 NAND2X1_396 ( .A(_1069_), .B(_1048_), .Y(_1072_) );
	OAI21X1 OAI21X1_793 ( .A(_1030_), .B(_1072_), .C(_1071_), .Y(_1073_) );
	XOR2X1 XOR2X1_27 ( .A(gen_nonce_synth_rand_20_), .B(_2__20_), .Y(_1074_) );
	NAND2X1 NAND2X1_397 ( .A(_1074_), .B(_1073_), .Y(_1075_) );
	OR2X2 OR2X2_31 ( .A(_1073_), .B(_1074_), .Y(_1076_) );
	AOI21X1 AOI21X1_616 ( .A(_1075_), .B(_1076_), .C(comparador_valid_bF_buf3), .Y(_1077_) );
	OAI21X1 OAI21X1_794 ( .A(_855__bF_buf1), .B(_2__20_), .C(_868__bF_buf2), .Y(_1078_) );
	OAI22X1 OAI22X1_225 ( .A(_854_), .B(_1066_), .C(_1077_), .D(_1078_), .Y(_827__20_) );
	INVX1 INVX1_643 ( .A(_2__21_), .Y(_1079_) );
	OAI21X1 OAI21X1_795 ( .A(_846_), .B(_1066_), .C(_1075_), .Y(_1080_) );
	NOR2X1 NOR2X1_256 ( .A(_847_), .B(_1079_), .Y(_1081_) );
	NOR2X1 NOR2X1_257 ( .A(gen_nonce_synth_rand_21_), .B(_2__21_), .Y(_1082_) );
	NOR2X1 NOR2X1_258 ( .A(_1082_), .B(_1081_), .Y(_1083_) );
	NAND2X1 NAND2X1_398 ( .A(_1083_), .B(_1080_), .Y(_1084_) );
	OR2X2 OR2X2_32 ( .A(_1080_), .B(_1083_), .Y(_1085_) );
	NAND3X1 NAND3X1_136 ( .A(_855__bF_buf0), .B(_1084_), .C(_1085_), .Y(_1086_) );
	AOI21X1 AOI21X1_617 ( .A(comparador_valid_bF_buf2), .B(_2__21_), .C(_867_), .Y(_1087_) );
	AOI22X1 AOI22X1_24 ( .A(_1__bF_buf3), .B(_1079_), .C(_1086_), .D(_1087_), .Y(_827__21_) );
	NAND2X1 NAND2X1_399 ( .A(_1__bF_buf2), .B(_2__22_), .Y(_1088_) );
	NAND2X1 NAND2X1_400 ( .A(gen_nonce_synth_rand_22_), .B(_2__22_), .Y(_1089_) );
	INVX1 INVX1_644 ( .A(_1089_), .Y(_1090_) );
	NOR2X1 NOR2X1_259 ( .A(gen_nonce_synth_rand_22_), .B(_2__22_), .Y(_1091_) );
	OR2X2 OR2X2_33 ( .A(_1090_), .B(_1091_), .Y(_1092_) );
	AND2X2 AND2X2_51 ( .A(_1083_), .B(_1074_), .Y(_1093_) );
	NAND2X1 NAND2X1_401 ( .A(_1093_), .B(_1073_), .Y(_1094_) );
	NAND2X1 NAND2X1_402 ( .A(gen_nonce_synth_rand_20_), .B(_2__20_), .Y(_1095_) );
	INVX1 INVX1_645 ( .A(_1081_), .Y(_1096_) );
	OAI21X1 OAI21X1_796 ( .A(_1082_), .B(_1095_), .C(_1096_), .Y(_1097_) );
	INVX1 INVX1_646 ( .A(_1097_), .Y(_1098_) );
	NAND3X1 NAND3X1_137 ( .A(_1092_), .B(_1098_), .C(_1094_), .Y(_1099_) );
	INVX1 INVX1_647 ( .A(_1092_), .Y(_1100_) );
	AND2X2 AND2X2_52 ( .A(_1073_), .B(_1093_), .Y(_1101_) );
	OAI21X1 OAI21X1_797 ( .A(_1101_), .B(_1097_), .C(_1100_), .Y(_1102_) );
	AOI21X1 AOI21X1_618 ( .A(_1099_), .B(_1102_), .C(comparador_valid_bF_buf1), .Y(_1103_) );
	OAI21X1 OAI21X1_798 ( .A(_855__bF_buf4), .B(_2__22_), .C(_868__bF_buf1), .Y(_1104_) );
	OAI21X1 OAI21X1_799 ( .A(_1103_), .B(_1104_), .C(_1088_), .Y(_827__22_) );
	INVX1 INVX1_648 ( .A(_2__23_), .Y(_1105_) );
	AOI21X1 AOI21X1_619 ( .A(_1098_), .B(_1094_), .C(_1092_), .Y(_1106_) );
	NOR2X1 NOR2X1_260 ( .A(_849_), .B(_1105_), .Y(_1107_) );
	NOR2X1 NOR2X1_261 ( .A(gen_nonce_synth_rand_23_), .B(_2__23_), .Y(_1108_) );
	OR2X2 OR2X2_34 ( .A(_1107_), .B(_1108_), .Y(_1109_) );
	INVX1 INVX1_649 ( .A(_1109_), .Y(_1110_) );
	OAI21X1 OAI21X1_800 ( .A(_1106_), .B(_1090_), .C(_1110_), .Y(_1111_) );
	NAND3X1 NAND3X1_138 ( .A(_1089_), .B(_1109_), .C(_1102_), .Y(_1112_) );
	NAND3X1 NAND3X1_139 ( .A(_855__bF_buf3), .B(_1111_), .C(_1112_), .Y(_1113_) );
	AOI21X1 AOI21X1_620 ( .A(comparador_valid_bF_buf0), .B(_2__23_), .C(_867_), .Y(_1114_) );
	AOI22X1 AOI22X1_25 ( .A(_1__bF_buf1), .B(_1105_), .C(_1113_), .D(_1114_), .Y(_827__23_) );
	INVX1 INVX1_650 ( .A(_2__24_), .Y(_1115_) );
	NAND2X1 NAND2X1_403 ( .A(gen_nonce_synth_rand_8_), .B(_933_), .Y(_1116_) );
	NAND2X1 NAND2X1_404 ( .A(_2__8_), .B(_834_), .Y(_1117_) );
	NAND2X1 NAND2X1_405 ( .A(gen_nonce_synth_rand_9_), .B(_947_), .Y(_1118_) );
	NAND2X1 NAND2X1_406 ( .A(_2__9_), .B(_835_), .Y(_1119_) );
	AOI22X1 AOI22X1_26 ( .A(_1116_), .B(_1117_), .C(_1118_), .D(_1119_), .Y(_1120_) );
	NAND3X1 NAND3X1_140 ( .A(_960_), .B(_969_), .C(_1120_), .Y(_1121_) );
	NOR3X1 NOR3X1_7 ( .A(_998_), .B(_1021_), .C(_1121_), .Y(_1122_) );
	NAND2X1 NAND2X1_407 ( .A(_941_), .B(_1122_), .Y(_1123_) );
	NOR2X1 NOR2X1_262 ( .A(_1092_), .B(_1109_), .Y(_1124_) );
	NAND2X1 NAND2X1_408 ( .A(_1093_), .B(_1124_), .Y(_1125_) );
	OR2X2 OR2X2_35 ( .A(_1072_), .B(_1125_), .Y(_1126_) );
	AOI21X1 AOI21X1_621 ( .A(_1028_), .B(_1123_), .C(_1126_), .Y(_1127_) );
	NOR2X1 NOR2X1_263 ( .A(_1071_), .B(_1125_), .Y(_1128_) );
	AOI21X1 AOI21X1_622 ( .A(_1090_), .B(_1110_), .C(_1107_), .Y(_1129_) );
	NAND2X1 NAND2X1_409 ( .A(_1097_), .B(_1124_), .Y(_1130_) );
	NAND2X1 NAND2X1_410 ( .A(_1129_), .B(_1130_), .Y(_1131_) );
	OR2X2 OR2X2_36 ( .A(_1128_), .B(_1131_), .Y(_1132_) );
	NOR2X1 NOR2X1_264 ( .A(_850_), .B(_1115_), .Y(_1133_) );
	INVX1 INVX1_651 ( .A(_1133_), .Y(_1134_) );
	NAND2X1 NAND2X1_411 ( .A(_850_), .B(_1115_), .Y(_1135_) );
	NAND2X1 NAND2X1_412 ( .A(_1135_), .B(_1134_), .Y(_1136_) );
	INVX1 INVX1_652 ( .A(_1136_), .Y(_1137_) );
	OAI21X1 OAI21X1_801 ( .A(_1127_), .B(_1132_), .C(_1137_), .Y(_1138_) );
	NOR2X1 NOR2X1_265 ( .A(_1132_), .B(_1127_), .Y(_1139_) );
	NAND2X1 NAND2X1_413 ( .A(_1136_), .B(_1139_), .Y(_1140_) );
	AOI21X1 AOI21X1_623 ( .A(_1138_), .B(_1140_), .C(comparador_valid_bF_buf5), .Y(_1141_) );
	OAI21X1 OAI21X1_802 ( .A(_855__bF_buf2), .B(_2__24_), .C(_868__bF_buf0), .Y(_1142_) );
	OAI22X1 OAI22X1_226 ( .A(_854_), .B(_1115_), .C(_1141_), .D(_1142_), .Y(_827__24_) );
	NAND2X1 NAND2X1_414 ( .A(_1__bF_buf0), .B(_2__25_), .Y(_1143_) );
	NAND2X1 NAND2X1_415 ( .A(gen_nonce_synth_rand_25_), .B(_2__25_), .Y(_1144_) );
	INVX1 INVX1_653 ( .A(_1144_), .Y(_1145_) );
	NOR2X1 NOR2X1_266 ( .A(gen_nonce_synth_rand_25_), .B(_2__25_), .Y(_1146_) );
	NOR2X1 NOR2X1_267 ( .A(_1146_), .B(_1145_), .Y(_1147_) );
	OAI21X1 OAI21X1_803 ( .A(_850_), .B(_1115_), .C(_1138_), .Y(_1148_) );
	OR2X2 OR2X2_37 ( .A(_1148_), .B(_1147_), .Y(_1149_) );
	INVX1 INVX1_654 ( .A(_1147_), .Y(_1150_) );
	NOR2X1 NOR2X1_268 ( .A(_1136_), .B(_1150_), .Y(_1151_) );
	OAI21X1 OAI21X1_804 ( .A(_1127_), .B(_1132_), .C(_1151_), .Y(_1152_) );
	OAI21X1 OAI21X1_805 ( .A(_1134_), .B(_1150_), .C(_1152_), .Y(_1153_) );
	INVX1 INVX1_655 ( .A(_1153_), .Y(_1154_) );
	AOI21X1 AOI21X1_624 ( .A(_1154_), .B(_1149_), .C(comparador_valid_bF_buf4), .Y(_1155_) );
	OAI21X1 OAI21X1_806 ( .A(_855__bF_buf1), .B(_2__25_), .C(_868__bF_buf3), .Y(_1156_) );
	OAI21X1 OAI21X1_807 ( .A(_1155_), .B(_1156_), .C(_1143_), .Y(_827__25_) );
	NAND2X1 NAND2X1_416 ( .A(_1__bF_buf5), .B(_2__26_), .Y(_1157_) );
	OAI21X1 OAI21X1_808 ( .A(_1134_), .B(_1146_), .C(_1144_), .Y(_1158_) );
	INVX1 INVX1_656 ( .A(_1158_), .Y(_1159_) );
	XNOR2X1 XNOR2X1_25 ( .A(gen_nonce_synth_rand_26_), .B(_2__26_), .Y(_1160_) );
	NAND3X1 NAND3X1_141 ( .A(_1159_), .B(_1160_), .C(_1152_), .Y(_1161_) );
	AOI21X1 AOI21X1_625 ( .A(_1159_), .B(_1152_), .C(_1160_), .Y(_1162_) );
	INVX1 INVX1_657 ( .A(_1162_), .Y(_1163_) );
	AOI21X1 AOI21X1_626 ( .A(_1161_), .B(_1163_), .C(comparador_valid_bF_buf3), .Y(_1164_) );
	OAI21X1 OAI21X1_809 ( .A(_855__bF_buf0), .B(_2__26_), .C(_868__bF_buf2), .Y(_1165_) );
	OAI21X1 OAI21X1_810 ( .A(_1164_), .B(_1165_), .C(_1157_), .Y(_827__26_) );
	NAND2X1 NAND2X1_417 ( .A(gen_nonce_synth_rand_26_), .B(_2__26_), .Y(_1166_) );
	INVX1 INVX1_658 ( .A(_1166_), .Y(_1167_) );
	NAND2X1 NAND2X1_418 ( .A(gen_nonce_synth_rand_27_), .B(_2__27_), .Y(_1168_) );
	INVX1 INVX1_659 ( .A(_1168_), .Y(_1169_) );
	NOR2X1 NOR2X1_269 ( .A(gen_nonce_synth_rand_27_), .B(_2__27_), .Y(_1170_) );
	NOR2X1 NOR2X1_270 ( .A(_1170_), .B(_1169_), .Y(_1171_) );
	OAI21X1 OAI21X1_811 ( .A(_1162_), .B(_1167_), .C(_1171_), .Y(_1172_) );
	NOR2X1 NOR2X1_271 ( .A(_1167_), .B(_1162_), .Y(_1173_) );
	OAI21X1 OAI21X1_812 ( .A(_1169_), .B(_1170_), .C(_1173_), .Y(_1174_) );
	AOI21X1 AOI21X1_627 ( .A(_1172_), .B(_1174_), .C(comparador_valid_bF_buf2), .Y(_1175_) );
	OAI21X1 OAI21X1_813 ( .A(_855__bF_buf4), .B(_2__27_), .C(_868__bF_buf1), .Y(_1176_) );
	NAND2X1 NAND2X1_419 ( .A(_1__bF_buf4), .B(_2__27_), .Y(_1177_) );
	OAI21X1 OAI21X1_814 ( .A(_1175_), .B(_1176_), .C(_1177_), .Y(_827__27_) );
	INVX1 INVX1_660 ( .A(_2__28_), .Y(_1178_) );
	INVX1 INVX1_661 ( .A(_1160_), .Y(_1179_) );
	NAND2X1 NAND2X1_420 ( .A(_1171_), .B(_1179_), .Y(_1180_) );
	INVX1 INVX1_662 ( .A(_1180_), .Y(_1181_) );
	NAND2X1 NAND2X1_421 ( .A(_1181_), .B(_1151_), .Y(_1182_) );
	OAI21X1 OAI21X1_815 ( .A(_1170_), .B(_1166_), .C(_1168_), .Y(_1183_) );
	INVX1 INVX1_663 ( .A(_1183_), .Y(_1184_) );
	OAI21X1 OAI21X1_816 ( .A(_1159_), .B(_1180_), .C(_1184_), .Y(_1185_) );
	INVX1 INVX1_664 ( .A(_1185_), .Y(_1186_) );
	OAI21X1 OAI21X1_817 ( .A(_1139_), .B(_1182_), .C(_1186_), .Y(_1187_) );
	NOR2X1 NOR2X1_272 ( .A(_852_), .B(_1178_), .Y(_1188_) );
	INVX1 INVX1_665 ( .A(_1188_), .Y(_1189_) );
	NAND2X1 NAND2X1_422 ( .A(_852_), .B(_1178_), .Y(_1190_) );
	AND2X2 AND2X2_53 ( .A(_1189_), .B(_1190_), .Y(_1191_) );
	NOR2X1 NOR2X1_273 ( .A(_1191_), .B(_1187_), .Y(_1192_) );
	NOR2X1 NOR2X1_274 ( .A(_1072_), .B(_1125_), .Y(_1193_) );
	OAI21X1 OAI21X1_818 ( .A(_1024_), .B(_1029_), .C(_1193_), .Y(_1194_) );
	NOR2X1 NOR2X1_275 ( .A(_1131_), .B(_1128_), .Y(_1195_) );
	AOI21X1 AOI21X1_628 ( .A(_1195_), .B(_1194_), .C(_1182_), .Y(_1196_) );
	OAI21X1 OAI21X1_819 ( .A(_1196_), .B(_1185_), .C(_1191_), .Y(_1197_) );
	INVX1 INVX1_666 ( .A(_1197_), .Y(_1198_) );
	OAI21X1 OAI21X1_820 ( .A(_1192_), .B(_1198_), .C(_855__bF_buf3), .Y(_1199_) );
	OAI21X1 OAI21X1_821 ( .A(_855__bF_buf2), .B(_2__28_), .C(_1199_), .Y(_1200_) );
	OAI22X1 OAI22X1_227 ( .A(_854_), .B(_1178_), .C(_1200_), .D(_867_), .Y(_827__28_) );
	INVX1 INVX1_667 ( .A(_2__29_), .Y(_1201_) );
	OAI21X1 OAI21X1_822 ( .A(_852_), .B(_1178_), .C(_1197_), .Y(_1202_) );
	NOR2X1 NOR2X1_276 ( .A(_853_), .B(_1201_), .Y(_1203_) );
	NOR2X1 NOR2X1_277 ( .A(gen_nonce_synth_rand_29_), .B(_2__29_), .Y(_1204_) );
	NOR2X1 NOR2X1_278 ( .A(_1204_), .B(_1203_), .Y(_1205_) );
	INVX1 INVX1_668 ( .A(_1205_), .Y(_1206_) );
	OAI21X1 OAI21X1_823 ( .A(_1202_), .B(_1206_), .C(_855__bF_buf1), .Y(_1207_) );
	AOI21X1 AOI21X1_629 ( .A(_1202_), .B(_1206_), .C(_1207_), .Y(_1208_) );
	OAI21X1 OAI21X1_824 ( .A(_855__bF_buf0), .B(_2__29_), .C(_868__bF_buf0), .Y(_1209_) );
	OAI22X1 OAI22X1_228 ( .A(_854_), .B(_1201_), .C(_1208_), .D(_1209_), .Y(_827__29_) );
	NAND2X1 NAND2X1_423 ( .A(_1__bF_buf3), .B(_2__30_), .Y(_1210_) );
	INVX1 INVX1_669 ( .A(_1182_), .Y(_1211_) );
	OAI21X1 OAI21X1_825 ( .A(_1127_), .B(_1132_), .C(_1211_), .Y(_1212_) );
	INVX1 INVX1_670 ( .A(_1191_), .Y(_1213_) );
	NOR2X1 NOR2X1_279 ( .A(_1206_), .B(_1213_), .Y(_1214_) );
	INVX1 INVX1_671 ( .A(_1214_), .Y(_1215_) );
	AOI21X1 AOI21X1_630 ( .A(_1186_), .B(_1212_), .C(_1215_), .Y(_1216_) );
	AOI21X1 AOI21X1_631 ( .A(_1188_), .B(_1205_), .C(_1203_), .Y(_1217_) );
	INVX1 INVX1_672 ( .A(_1217_), .Y(_1218_) );
	NAND2X1 NAND2X1_424 ( .A(gen_nonce_synth_rand_30_), .B(_2__30_), .Y(_1219_) );
	INVX1 INVX1_673 ( .A(_1219_), .Y(_1220_) );
	NOR2X1 NOR2X1_280 ( .A(gen_nonce_synth_rand_30_), .B(_2__30_), .Y(_1221_) );
	NOR2X1 NOR2X1_281 ( .A(_1221_), .B(_1220_), .Y(_1222_) );
	OAI21X1 OAI21X1_826 ( .A(_1216_), .B(_1218_), .C(_1222_), .Y(_1223_) );
	OAI21X1 OAI21X1_827 ( .A(_1196_), .B(_1185_), .C(_1214_), .Y(_1224_) );
	INVX1 INVX1_674 ( .A(_1222_), .Y(_1225_) );
	NAND3X1 NAND3X1_142 ( .A(_1217_), .B(_1225_), .C(_1224_), .Y(_1226_) );
	AOI21X1 AOI21X1_632 ( .A(_1226_), .B(_1223_), .C(comparador_valid_bF_buf1), .Y(_1227_) );
	OAI21X1 OAI21X1_828 ( .A(_855__bF_buf4), .B(_2__30_), .C(_868__bF_buf3), .Y(_1228_) );
	OAI21X1 OAI21X1_829 ( .A(_1227_), .B(_1228_), .C(_1210_), .Y(_827__30_) );
	AOI21X1 AOI21X1_633 ( .A(_1217_), .B(_1224_), .C(_1225_), .Y(_1229_) );
	XNOR2X1 XNOR2X1_26 ( .A(gen_nonce_synth_rand_31_), .B(_2__31_), .Y(_1230_) );
	INVX1 INVX1_675 ( .A(_1230_), .Y(_1231_) );
	OAI21X1 OAI21X1_830 ( .A(_1229_), .B(_1220_), .C(_1231_), .Y(_1232_) );
	NAND3X1 NAND3X1_143 ( .A(_1219_), .B(_1230_), .C(_1223_), .Y(_1233_) );
	NAND3X1 NAND3X1_144 ( .A(_855__bF_buf3), .B(_1233_), .C(_1232_), .Y(_1234_) );
	AOI21X1 AOI21X1_634 ( .A(comparador_valid_bF_buf0), .B(_2__31_), .C(_867_), .Y(_1235_) );
	NOR2X1 NOR2X1_282 ( .A(_2__31_), .B(_854_), .Y(_1236_) );
	AOI21X1 AOI21X1_635 ( .A(_1235_), .B(_1234_), .C(_1236_), .Y(_827__31_) );
	DFFPOSX1 DFFPOSX1_815 ( .CLK(clk_bF_buf97), .D(_827__0_), .Q(_2__0_) );
	DFFPOSX1 DFFPOSX1_816 ( .CLK(clk_bF_buf96), .D(_827__1_), .Q(_2__1_) );
	DFFPOSX1 DFFPOSX1_817 ( .CLK(clk_bF_buf95), .D(_827__2_), .Q(_2__2_) );
	DFFPOSX1 DFFPOSX1_818 ( .CLK(clk_bF_buf94), .D(_827__3_), .Q(_2__3_) );
	DFFPOSX1 DFFPOSX1_819 ( .CLK(clk_bF_buf93), .D(_827__4_), .Q(_2__4_) );
	DFFPOSX1 DFFPOSX1_820 ( .CLK(clk_bF_buf92), .D(_827__5_), .Q(_2__5_) );
	DFFPOSX1 DFFPOSX1_821 ( .CLK(clk_bF_buf91), .D(_827__6_), .Q(_2__6_) );
	DFFPOSX1 DFFPOSX1_822 ( .CLK(clk_bF_buf90), .D(_827__7_), .Q(_2__7_) );
	DFFPOSX1 DFFPOSX1_823 ( .CLK(clk_bF_buf89), .D(_827__8_), .Q(_2__8_) );
	DFFPOSX1 DFFPOSX1_824 ( .CLK(clk_bF_buf88), .D(_827__9_), .Q(_2__9_) );
	DFFPOSX1 DFFPOSX1_825 ( .CLK(clk_bF_buf87), .D(_827__10_), .Q(_2__10_) );
	DFFPOSX1 DFFPOSX1_826 ( .CLK(clk_bF_buf86), .D(_827__11_), .Q(_2__11_) );
	DFFPOSX1 DFFPOSX1_827 ( .CLK(clk_bF_buf85), .D(_827__12_), .Q(_2__12_) );
	DFFPOSX1 DFFPOSX1_828 ( .CLK(clk_bF_buf84), .D(_827__13_), .Q(_2__13_) );
	DFFPOSX1 DFFPOSX1_829 ( .CLK(clk_bF_buf83), .D(_827__14_), .Q(_2__14_) );
	DFFPOSX1 DFFPOSX1_830 ( .CLK(clk_bF_buf82), .D(_827__15_), .Q(_2__15_) );
	DFFPOSX1 DFFPOSX1_831 ( .CLK(clk_bF_buf81), .D(_827__16_), .Q(_2__16_) );
	DFFPOSX1 DFFPOSX1_832 ( .CLK(clk_bF_buf80), .D(_827__17_), .Q(_2__17_) );
	DFFPOSX1 DFFPOSX1_833 ( .CLK(clk_bF_buf79), .D(_827__18_), .Q(_2__18_) );
	DFFPOSX1 DFFPOSX1_834 ( .CLK(clk_bF_buf78), .D(_827__19_), .Q(_2__19_) );
	DFFPOSX1 DFFPOSX1_835 ( .CLK(clk_bF_buf77), .D(_827__20_), .Q(_2__20_) );
	DFFPOSX1 DFFPOSX1_836 ( .CLK(clk_bF_buf76), .D(_827__21_), .Q(_2__21_) );
	DFFPOSX1 DFFPOSX1_837 ( .CLK(clk_bF_buf75), .D(_827__22_), .Q(_2__22_) );
	DFFPOSX1 DFFPOSX1_838 ( .CLK(clk_bF_buf74), .D(_827__23_), .Q(_2__23_) );
	DFFPOSX1 DFFPOSX1_839 ( .CLK(clk_bF_buf73), .D(_827__24_), .Q(_2__24_) );
	DFFPOSX1 DFFPOSX1_840 ( .CLK(clk_bF_buf72), .D(_827__25_), .Q(_2__25_) );
	DFFPOSX1 DFFPOSX1_841 ( .CLK(clk_bF_buf71), .D(_827__26_), .Q(_2__26_) );
	DFFPOSX1 DFFPOSX1_842 ( .CLK(clk_bF_buf70), .D(_827__27_), .Q(_2__27_) );
	DFFPOSX1 DFFPOSX1_843 ( .CLK(clk_bF_buf69), .D(_827__28_), .Q(_2__28_) );
	DFFPOSX1 DFFPOSX1_844 ( .CLK(clk_bF_buf68), .D(_827__29_), .Q(_2__29_) );
	DFFPOSX1 DFFPOSX1_845 ( .CLK(clk_bF_buf67), .D(_827__30_), .Q(_2__30_) );
	DFFPOSX1 DFFPOSX1_846 ( .CLK(clk_bF_buf66), .D(_827__31_), .Q(_2__31_) );
	DFFPOSX1 DFFPOSX1_847 ( .CLK(clk_bF_buf65), .D(_828__0_), .Q(gen_nonce_synth_rand_0_) );
	DFFPOSX1 DFFPOSX1_848 ( .CLK(clk_bF_buf64), .D(_828__1_), .Q(gen_nonce_synth_rand_1_) );
	DFFPOSX1 DFFPOSX1_849 ( .CLK(clk_bF_buf63), .D(_828__2_), .Q(gen_nonce_synth_rand_2_) );
	DFFPOSX1 DFFPOSX1_850 ( .CLK(clk_bF_buf62), .D(_828__3_), .Q(gen_nonce_synth_rand_3_) );
	DFFPOSX1 DFFPOSX1_851 ( .CLK(clk_bF_buf61), .D(_828__4_), .Q(gen_nonce_synth_rand_4_) );
	DFFPOSX1 DFFPOSX1_852 ( .CLK(clk_bF_buf60), .D(_828__5_), .Q(gen_nonce_synth_rand_5_) );
	DFFPOSX1 DFFPOSX1_853 ( .CLK(clk_bF_buf59), .D(_828__6_), .Q(gen_nonce_synth_rand_6_) );
	DFFPOSX1 DFFPOSX1_854 ( .CLK(clk_bF_buf58), .D(_828__7_), .Q(gen_nonce_synth_rand_7_) );
	DFFPOSX1 DFFPOSX1_855 ( .CLK(clk_bF_buf57), .D(_828__8_), .Q(gen_nonce_synth_rand_8_) );
	DFFPOSX1 DFFPOSX1_856 ( .CLK(clk_bF_buf56), .D(_828__9_), .Q(gen_nonce_synth_rand_9_) );
	DFFPOSX1 DFFPOSX1_857 ( .CLK(clk_bF_buf55), .D(_828__10_), .Q(gen_nonce_synth_rand_10_) );
	DFFPOSX1 DFFPOSX1_858 ( .CLK(clk_bF_buf54), .D(_828__11_), .Q(gen_nonce_synth_rand_11_) );
	DFFPOSX1 DFFPOSX1_859 ( .CLK(clk_bF_buf53), .D(_828__12_), .Q(gen_nonce_synth_rand_12_) );
	DFFPOSX1 DFFPOSX1_860 ( .CLK(clk_bF_buf52), .D(_828__13_), .Q(gen_nonce_synth_rand_13_) );
	DFFPOSX1 DFFPOSX1_861 ( .CLK(clk_bF_buf51), .D(_828__14_), .Q(gen_nonce_synth_rand_14_) );
	DFFPOSX1 DFFPOSX1_862 ( .CLK(clk_bF_buf50), .D(_828__15_), .Q(gen_nonce_synth_rand_15_) );
	DFFPOSX1 DFFPOSX1_863 ( .CLK(clk_bF_buf49), .D(_828__16_), .Q(gen_nonce_synth_rand_16_) );
	DFFPOSX1 DFFPOSX1_864 ( .CLK(clk_bF_buf48), .D(_828__17_), .Q(gen_nonce_synth_rand_17_) );
	DFFPOSX1 DFFPOSX1_865 ( .CLK(clk_bF_buf47), .D(_828__18_), .Q(gen_nonce_synth_rand_18_) );
	DFFPOSX1 DFFPOSX1_866 ( .CLK(clk_bF_buf46), .D(_828__19_), .Q(gen_nonce_synth_rand_19_) );
	DFFPOSX1 DFFPOSX1_867 ( .CLK(clk_bF_buf45), .D(_828__20_), .Q(gen_nonce_synth_rand_20_) );
	DFFPOSX1 DFFPOSX1_868 ( .CLK(clk_bF_buf44), .D(_828__21_), .Q(gen_nonce_synth_rand_21_) );
	DFFPOSX1 DFFPOSX1_869 ( .CLK(clk_bF_buf43), .D(_828__22_), .Q(gen_nonce_synth_rand_22_) );
	DFFPOSX1 DFFPOSX1_870 ( .CLK(clk_bF_buf42), .D(_828__23_), .Q(gen_nonce_synth_rand_23_) );
	DFFPOSX1 DFFPOSX1_871 ( .CLK(clk_bF_buf41), .D(_828__24_), .Q(gen_nonce_synth_rand_24_) );
	DFFPOSX1 DFFPOSX1_872 ( .CLK(clk_bF_buf40), .D(_828__25_), .Q(gen_nonce_synth_rand_25_) );
	DFFPOSX1 DFFPOSX1_873 ( .CLK(clk_bF_buf39), .D(_828__26_), .Q(gen_nonce_synth_rand_26_) );
	DFFPOSX1 DFFPOSX1_874 ( .CLK(clk_bF_buf38), .D(_828__27_), .Q(gen_nonce_synth_rand_27_) );
	DFFPOSX1 DFFPOSX1_875 ( .CLK(clk_bF_buf37), .D(_828__28_), .Q(gen_nonce_synth_rand_28_) );
	DFFPOSX1 DFFPOSX1_876 ( .CLK(clk_bF_buf36), .D(_828__29_), .Q(gen_nonce_synth_rand_29_) );
	DFFPOSX1 DFFPOSX1_877 ( .CLK(clk_bF_buf35), .D(_828__30_), .Q(gen_nonce_synth_rand_30_) );
	DFFPOSX1 DFFPOSX1_878 ( .CLK(clk_bF_buf34), .D(_828__31_), .Q(gen_nonce_synth_rand_31_) );
	INVX1 INVX1_676 ( .A(micro_hash_synth_1_W_26__0_), .Y(_2918_) );
	OR2X2 OR2X2_38 ( .A(concatenador_counter_3_), .B(concatenador_counter_2_), .Y(_2919_) );
	NOR2X1 NOR2X1_283 ( .A(concatenador_counter_5_), .B(concatenador_counter_4_), .Y(_2920_) );
	INVX1 INVX1_677 ( .A(_2920_), .Y(_2921_) );
	NOR2X1 NOR2X1_284 ( .A(_2919_), .B(_2921_), .Y(_2922_) );
	INVX8 INVX8_6 ( .A(concatenador_counter_0_bF_buf1), .Y(_2923_) );
	NOR2X1 NOR2X1_285 ( .A(concatenador_counter_1_bF_buf5), .B(_2923__bF_buf7), .Y(_2924_) );
	NAND3X1 NAND3X1_145 ( .A(reset_L_bF_buf6), .B(_2924_), .C(_2922_), .Y(_2925_) );
	NOR2X1 NOR2X1_286 ( .A(concatenador_counter_1_bF_buf4), .B(_2919_), .Y(_2926_) );
	INVX1 INVX1_678 ( .A(_2926_), .Y(_2927_) );
	NOR2X1 NOR2X1_287 ( .A(_2921_), .B(_2927_), .Y(_2928_) );
	INVX1 INVX1_679 ( .A(_2928_), .Y(_2929_) );
	OAI21X1 OAI21X1_831 ( .A(_2929_), .B(_2923__bF_buf6), .C(reset_L_bF_buf5), .Y(_2930_) );
	XOR2X1 XOR2X1_28 ( .A(micro_hash_synth_1_W_12__0_), .B(micro_hash_synth_1_W_17__0_), .Y(_2931_) );
	NOR2X1 NOR2X1_288 ( .A(micro_hash_synth_1_W_23__0_), .B(_2931_), .Y(_2932_) );
	OAI22X1 OAI22X1_229 ( .A(_2925__bF_buf15), .B(_2932_), .C(_2930__bF_buf13), .D(_2918_), .Y(_1400_) );
	INVX1 INVX1_680 ( .A(micro_hash_synth_1_W_26__1_), .Y(_2933_) );
	INVX1 INVX1_681 ( .A(micro_hash_synth_1_W_12__1_), .Y(_2934_) );
	INVX1 INVX1_682 ( .A(micro_hash_synth_1_W_23__1_), .Y(_2935_) );
	OAI21X1 OAI21X1_832 ( .A(_2934_), .B(micro_hash_synth_1_W_17__1_), .C(_2935_), .Y(_2936_) );
	AOI21X1 AOI21X1_636 ( .A(_2934_), .B(micro_hash_synth_1_W_17__1_), .C(_2936_), .Y(_2937_) );
	OAI22X1 OAI22X1_230 ( .A(_2925__bF_buf14), .B(_2937_), .C(_2930__bF_buf12), .D(_2933_), .Y(_1401_) );
	INVX1 INVX1_683 ( .A(micro_hash_synth_1_W_26__2_), .Y(_2938_) );
	INVX1 INVX1_684 ( .A(micro_hash_synth_1_W_12__2_), .Y(_2939_) );
	INVX1 INVX1_685 ( .A(micro_hash_synth_1_W_23__2_), .Y(_2940_) );
	OAI21X1 OAI21X1_833 ( .A(_2939_), .B(micro_hash_synth_1_W_17__2_), .C(_2940_), .Y(_2941_) );
	AOI21X1 AOI21X1_637 ( .A(_2939_), .B(micro_hash_synth_1_W_17__2_), .C(_2941_), .Y(_2942_) );
	OAI22X1 OAI22X1_231 ( .A(_2925__bF_buf13), .B(_2942_), .C(_2930__bF_buf11), .D(_2938_), .Y(_1402_) );
	INVX1 INVX1_686 ( .A(micro_hash_synth_1_W_26__3_), .Y(_2943_) );
	XOR2X1 XOR2X1_29 ( .A(micro_hash_synth_1_W_12__3_), .B(micro_hash_synth_1_W_17__3_), .Y(_2944_) );
	NOR2X1 NOR2X1_289 ( .A(micro_hash_synth_1_W_23__3_), .B(_2944_), .Y(_2945_) );
	OAI22X1 OAI22X1_232 ( .A(_2925__bF_buf12), .B(_2945_), .C(_2930__bF_buf10), .D(_2943_), .Y(_1403_) );
	INVX1 INVX1_687 ( .A(micro_hash_synth_1_W_26__4_), .Y(_2946_) );
	XOR2X1 XOR2X1_30 ( .A(micro_hash_synth_1_W_12__4_), .B(micro_hash_synth_1_W_17__4_), .Y(_2947_) );
	NOR2X1 NOR2X1_290 ( .A(micro_hash_synth_1_W_23__4_), .B(_2947_), .Y(_2948_) );
	OAI22X1 OAI22X1_233 ( .A(_2925__bF_buf11), .B(_2948_), .C(_2930__bF_buf9), .D(_2946_), .Y(_1404_) );
	INVX1 INVX1_688 ( .A(micro_hash_synth_1_W_26__5_), .Y(_2949_) );
	XOR2X1 XOR2X1_31 ( .A(micro_hash_synth_1_W_12__5_), .B(micro_hash_synth_1_W_17__5_), .Y(_2950_) );
	NOR2X1 NOR2X1_291 ( .A(micro_hash_synth_1_W_23__5_), .B(_2950_), .Y(_2951_) );
	OAI22X1 OAI22X1_234 ( .A(_2925__bF_buf10), .B(_2951_), .C(_2930__bF_buf8), .D(_2949_), .Y(_1405_) );
	INVX1 INVX1_689 ( .A(micro_hash_synth_1_W_26__6_), .Y(_2952_) );
	INVX1 INVX1_690 ( .A(micro_hash_synth_1_W_12__6_), .Y(_2953_) );
	INVX1 INVX1_691 ( .A(micro_hash_synth_1_W_23__6_), .Y(_2954_) );
	OAI21X1 OAI21X1_834 ( .A(_2953_), .B(micro_hash_synth_1_W_17__6_), .C(_2954_), .Y(_2955_) );
	AOI21X1 AOI21X1_638 ( .A(_2953_), .B(micro_hash_synth_1_W_17__6_), .C(_2955_), .Y(_2956_) );
	OAI22X1 OAI22X1_235 ( .A(_2925__bF_buf9), .B(_2956_), .C(_2930__bF_buf7), .D(_2952_), .Y(_1412_) );
	INVX1 INVX1_692 ( .A(micro_hash_synth_1_W_26__7_), .Y(_2957_) );
	INVX1 INVX1_693 ( .A(micro_hash_synth_1_W_12__7_), .Y(_2958_) );
	INVX1 INVX1_694 ( .A(micro_hash_synth_1_W_23__7_), .Y(_2959_) );
	OAI21X1 OAI21X1_835 ( .A(_2958_), .B(micro_hash_synth_1_W_17__7_), .C(_2959_), .Y(_2960_) );
	AOI21X1 AOI21X1_639 ( .A(_2958_), .B(micro_hash_synth_1_W_17__7_), .C(_2960_), .Y(_2961_) );
	OAI22X1 OAI22X1_236 ( .A(_2925__bF_buf8), .B(_2961_), .C(_2930__bF_buf6), .D(_2957_), .Y(_1423_) );
	INVX1 INVX1_695 ( .A(micro_hash_synth_1_W_25__0_), .Y(_2962_) );
	XOR2X1 XOR2X1_32 ( .A(micro_hash_synth_1_W_11__0_), .B(micro_hash_synth_1_W_16__0_), .Y(_2963_) );
	NOR2X1 NOR2X1_292 ( .A(micro_hash_synth_1_W_22__0_), .B(_2963_), .Y(_2964_) );
	OAI22X1 OAI22X1_237 ( .A(_2925__bF_buf7), .B(_2964_), .C(_2930__bF_buf5), .D(_2962_), .Y(_1434_) );
	INVX1 INVX1_696 ( .A(micro_hash_synth_1_W_25__1_), .Y(_2965_) );
	INVX1 INVX1_697 ( .A(micro_hash_synth_1_W_11__1_), .Y(_2966_) );
	INVX1 INVX1_698 ( .A(micro_hash_synth_1_W_22__1_), .Y(_2967_) );
	OAI21X1 OAI21X1_836 ( .A(_2966_), .B(micro_hash_synth_1_W_16__1_), .C(_2967_), .Y(_2968_) );
	AOI21X1 AOI21X1_640 ( .A(_2966_), .B(micro_hash_synth_1_W_16__1_), .C(_2968_), .Y(_2969_) );
	OAI22X1 OAI22X1_238 ( .A(_2925__bF_buf6), .B(_2969_), .C(_2930__bF_buf4), .D(_2965_), .Y(_1445_) );
	INVX1 INVX1_699 ( .A(micro_hash_synth_1_W_25__2_), .Y(_2970_) );
	INVX1 INVX1_700 ( .A(micro_hash_synth_1_W_11__2_), .Y(_2971_) );
	INVX1 INVX1_701 ( .A(micro_hash_synth_1_W_22__2_), .Y(_2972_) );
	OAI21X1 OAI21X1_837 ( .A(_2971_), .B(micro_hash_synth_1_W_16__2_), .C(_2972_), .Y(_2973_) );
	AOI21X1 AOI21X1_641 ( .A(_2971_), .B(micro_hash_synth_1_W_16__2_), .C(_2973_), .Y(_2974_) );
	OAI22X1 OAI22X1_239 ( .A(_2925__bF_buf5), .B(_2974_), .C(_2930__bF_buf3), .D(_2970_), .Y(_1456_) );
	INVX1 INVX1_702 ( .A(micro_hash_synth_1_W_25__3_), .Y(_2975_) );
	XOR2X1 XOR2X1_33 ( .A(micro_hash_synth_1_W_11__3_), .B(micro_hash_synth_1_W_16__3_), .Y(_2976_) );
	NOR2X1 NOR2X1_293 ( .A(micro_hash_synth_1_W_22__3_), .B(_2976_), .Y(_2977_) );
	OAI22X1 OAI22X1_240 ( .A(_2925__bF_buf4), .B(_2977_), .C(_2930__bF_buf2), .D(_2975_), .Y(_1467_) );
	INVX1 INVX1_703 ( .A(micro_hash_synth_1_W_25__4_), .Y(_2978_) );
	XOR2X1 XOR2X1_34 ( .A(micro_hash_synth_1_W_11__4_), .B(micro_hash_synth_1_W_16__4_), .Y(_2979_) );
	NOR2X1 NOR2X1_294 ( .A(micro_hash_synth_1_W_22__4_), .B(_2979_), .Y(_2980_) );
	OAI22X1 OAI22X1_241 ( .A(_2925__bF_buf3), .B(_2980_), .C(_2930__bF_buf1), .D(_2978_), .Y(_1478_) );
	INVX1 INVX1_704 ( .A(micro_hash_synth_1_W_25__5_), .Y(_2981_) );
	XOR2X1 XOR2X1_35 ( .A(micro_hash_synth_1_W_11__5_), .B(micro_hash_synth_1_W_16__5_), .Y(_2982_) );
	NOR2X1 NOR2X1_295 ( .A(micro_hash_synth_1_W_22__5_), .B(_2982_), .Y(_2983_) );
	OAI22X1 OAI22X1_242 ( .A(_2925__bF_buf2), .B(_2983_), .C(_2930__bF_buf0), .D(_2981_), .Y(_1485_) );
	INVX1 INVX1_705 ( .A(micro_hash_synth_1_W_25__6_), .Y(_2984_) );
	XOR2X1 XOR2X1_36 ( .A(micro_hash_synth_1_W_11__6_), .B(micro_hash_synth_1_W_16__6_), .Y(_2985_) );
	NOR2X1 NOR2X1_296 ( .A(micro_hash_synth_1_W_22__6_), .B(_2985_), .Y(_2986_) );
	OAI22X1 OAI22X1_243 ( .A(_2925__bF_buf1), .B(_2986_), .C(_2930__bF_buf13), .D(_2984_), .Y(_1486_) );
	INVX1 INVX1_706 ( .A(micro_hash_synth_1_W_25__7_), .Y(_2987_) );
	XOR2X1 XOR2X1_37 ( .A(micro_hash_synth_1_W_11__7_), .B(micro_hash_synth_1_W_16__7_), .Y(_2988_) );
	NOR2X1 NOR2X1_297 ( .A(micro_hash_synth_1_W_22__7_), .B(_2988_), .Y(_2989_) );
	OAI22X1 OAI22X1_244 ( .A(_2925__bF_buf0), .B(_2989_), .C(_2930__bF_buf12), .D(_2987_), .Y(_1487_) );
	INVX1 INVX1_707 ( .A(micro_hash_synth_1_W_8__0_), .Y(_2990_) );
	INVX1 INVX1_708 ( .A(bloque_in_64_), .Y(_2991_) );
	OAI22X1 OAI22X1_245 ( .A(_2991_), .B(_2925__bF_buf15), .C(_2930__bF_buf11), .D(_2990_), .Y(_1492_) );
	INVX1 INVX1_709 ( .A(micro_hash_synth_1_W_8__1_), .Y(_2992_) );
	INVX1 INVX1_710 ( .A(bloque_in_65_), .Y(_2993_) );
	OAI22X1 OAI22X1_246 ( .A(_2993_), .B(_2925__bF_buf14), .C(_2930__bF_buf10), .D(_2992_), .Y(_1497_) );
	INVX1 INVX1_711 ( .A(micro_hash_synth_1_W_8__2_), .Y(_2994_) );
	INVX1 INVX1_712 ( .A(bloque_in_66_), .Y(_2995_) );
	OAI22X1 OAI22X1_247 ( .A(_2995_), .B(_2925__bF_buf13), .C(_2930__bF_buf9), .D(_2994_), .Y(_1498_) );
	INVX1 INVX1_713 ( .A(micro_hash_synth_1_W_8__3_), .Y(_2996_) );
	INVX1 INVX1_714 ( .A(bloque_in_67_), .Y(_2997_) );
	OAI22X1 OAI22X1_248 ( .A(_2997_), .B(_2925__bF_buf12), .C(_2930__bF_buf8), .D(_2996_), .Y(_1499_) );
	INVX1 INVX1_715 ( .A(micro_hash_synth_1_W_8__4_), .Y(_2998_) );
	INVX1 INVX1_716 ( .A(bloque_in_68_), .Y(_2999_) );
	OAI22X1 OAI22X1_249 ( .A(_2999_), .B(_2925__bF_buf11), .C(_2930__bF_buf7), .D(_2998_), .Y(_1244_) );
	INVX1 INVX1_717 ( .A(micro_hash_synth_1_W_8__5_), .Y(_3000_) );
	INVX1 INVX1_718 ( .A(bloque_in_69_), .Y(_3001_) );
	OAI22X1 OAI22X1_250 ( .A(_3001_), .B(_2925__bF_buf10), .C(_2930__bF_buf6), .D(_3000_), .Y(_1245_) );
	INVX1 INVX1_719 ( .A(micro_hash_synth_1_W_8__6_), .Y(_3002_) );
	INVX1 INVX1_720 ( .A(bloque_in_70_), .Y(_3003_) );
	OAI22X1 OAI22X1_251 ( .A(_3003_), .B(_2925__bF_buf9), .C(_2930__bF_buf5), .D(_3002_), .Y(_1253_) );
	INVX1 INVX1_721 ( .A(micro_hash_synth_1_W_8__7_), .Y(_3004_) );
	INVX1 INVX1_722 ( .A(bloque_in_71_), .Y(_3005_) );
	OAI22X1 OAI22X1_252 ( .A(_3005_), .B(_2925__bF_buf8), .C(_2930__bF_buf4), .D(_3004_), .Y(_1255_) );
	INVX1 INVX1_723 ( .A(micro_hash_synth_1_W_3__0_), .Y(_3006_) );
	INVX1 INVX1_724 ( .A(bloque_in_24_), .Y(_3007_) );
	OAI22X1 OAI22X1_253 ( .A(_3007_), .B(_2925__bF_buf7), .C(_2930__bF_buf3), .D(_3006_), .Y(_1256_) );
	INVX1 INVX1_725 ( .A(micro_hash_synth_1_W_3__1_), .Y(_3008_) );
	INVX1 INVX1_726 ( .A(bloque_in_25_), .Y(_3009_) );
	OAI22X1 OAI22X1_254 ( .A(_3009_), .B(_2925__bF_buf6), .C(_2930__bF_buf2), .D(_3008_), .Y(_1257_) );
	INVX1 INVX1_727 ( .A(micro_hash_synth_1_W_3__2_), .Y(_3010_) );
	INVX1 INVX1_728 ( .A(bloque_in_26_), .Y(_3011_) );
	OAI22X1 OAI22X1_255 ( .A(_3011_), .B(_2925__bF_buf5), .C(_2930__bF_buf1), .D(_3010_), .Y(_1266_) );
	INVX1 INVX1_729 ( .A(micro_hash_synth_1_W_3__3_), .Y(_3012_) );
	INVX1 INVX1_730 ( .A(bloque_in_27_), .Y(_3013_) );
	OAI22X1 OAI22X1_256 ( .A(_3013_), .B(_2925__bF_buf4), .C(_2930__bF_buf0), .D(_3012_), .Y(_1269_) );
	INVX1 INVX1_731 ( .A(micro_hash_synth_1_W_3__4_), .Y(_3014_) );
	INVX1 INVX1_732 ( .A(bloque_in_28_), .Y(_3015_) );
	OAI22X1 OAI22X1_257 ( .A(_3015_), .B(_2925__bF_buf3), .C(_2930__bF_buf13), .D(_3014_), .Y(_1285_) );
	INVX1 INVX1_733 ( .A(micro_hash_synth_1_W_3__5_), .Y(_3016_) );
	INVX1 INVX1_734 ( .A(bloque_in_29_), .Y(_3017_) );
	OAI22X1 OAI22X1_258 ( .A(_3017_), .B(_2925__bF_buf2), .C(_2930__bF_buf12), .D(_3016_), .Y(_1301_) );
	INVX1 INVX1_735 ( .A(micro_hash_synth_1_W_3__6_), .Y(_3018_) );
	INVX1 INVX1_736 ( .A(bloque_in_30_), .Y(_3019_) );
	OAI22X1 OAI22X1_259 ( .A(_3019_), .B(_2925__bF_buf1), .C(_2930__bF_buf11), .D(_3018_), .Y(_1317_) );
	INVX1 INVX1_737 ( .A(micro_hash_synth_1_W_3__7_), .Y(_3020_) );
	INVX1 INVX1_738 ( .A(bloque_in_31_), .Y(_3021_) );
	OAI22X1 OAI22X1_260 ( .A(_3021_), .B(_2925__bF_buf0), .C(_2930__bF_buf10), .D(_3020_), .Y(_1333_) );
	INVX8 INVX8_7 ( .A(reset_L_bF_buf4), .Y(_3022_) );
	INVX1 INVX1_739 ( .A(micro_hash_synth_1_W_1__0_), .Y(_3023_) );
	NOR2X1 NOR2X1_298 ( .A(_3022__bF_buf5), .B(_3023_), .Y(_1242__8_) );
	INVX1 INVX1_740 ( .A(micro_hash_synth_1_W_1__1_), .Y(_3024_) );
	NOR2X1 NOR2X1_299 ( .A(_3022__bF_buf4), .B(_3024_), .Y(_1242__9_) );
	INVX1 INVX1_741 ( .A(micro_hash_synth_1_W_1__2_), .Y(_3025_) );
	NOR2X1 NOR2X1_300 ( .A(_3022__bF_buf3), .B(_3025_), .Y(_1242__10_) );
	INVX1 INVX1_742 ( .A(micro_hash_synth_1_W_1__3_), .Y(_3026_) );
	NOR2X1 NOR2X1_301 ( .A(_3022__bF_buf2), .B(_3026_), .Y(_1242__11_) );
	INVX1 INVX1_743 ( .A(micro_hash_synth_1_W_1__4_), .Y(_3027_) );
	NOR2X1 NOR2X1_302 ( .A(_3022__bF_buf1), .B(_3027_), .Y(_1242__12_) );
	INVX1 INVX1_744 ( .A(micro_hash_synth_1_W_1__5_), .Y(_3028_) );
	NOR2X1 NOR2X1_303 ( .A(_3022__bF_buf0), .B(_3028_), .Y(_1242__13_) );
	INVX1 INVX1_745 ( .A(micro_hash_synth_1_W_1__6_), .Y(_3029_) );
	NOR2X1 NOR2X1_304 ( .A(_3022__bF_buf5), .B(_3029_), .Y(_1242__14_) );
	INVX1 INVX1_746 ( .A(micro_hash_synth_1_W_1__7_), .Y(_3030_) );
	NOR2X1 NOR2X1_305 ( .A(_3022__bF_buf4), .B(_3030_), .Y(_1242__15_) );
	INVX1 INVX1_747 ( .A(micro_hash_synth_1_W_0__0_), .Y(_3031_) );
	NOR2X1 NOR2X1_306 ( .A(_3022__bF_buf3), .B(_3031_), .Y(_1242__0_) );
	INVX1 INVX1_748 ( .A(micro_hash_synth_1_W_0__1_), .Y(_3032_) );
	NOR2X1 NOR2X1_307 ( .A(_3022__bF_buf2), .B(_3032_), .Y(_1242__1_) );
	INVX1 INVX1_749 ( .A(micro_hash_synth_1_W_0__2_), .Y(_3033_) );
	NOR2X1 NOR2X1_308 ( .A(_3022__bF_buf1), .B(_3033_), .Y(_1242__2_) );
	INVX1 INVX1_750 ( .A(micro_hash_synth_1_W_0__3_), .Y(_3034_) );
	NOR2X1 NOR2X1_309 ( .A(_3022__bF_buf0), .B(_3034_), .Y(_1242__3_) );
	INVX1 INVX1_751 ( .A(micro_hash_synth_1_W_0__4_), .Y(_3035_) );
	NOR2X1 NOR2X1_310 ( .A(_3022__bF_buf5), .B(_3035_), .Y(_1242__4_) );
	INVX1 INVX1_752 ( .A(micro_hash_synth_1_W_0__5_), .Y(_3036_) );
	NOR2X1 NOR2X1_311 ( .A(_3022__bF_buf4), .B(_3036_), .Y(_1242__5_) );
	INVX1 INVX1_753 ( .A(micro_hash_synth_1_W_0__6_), .Y(_3037_) );
	NOR2X1 NOR2X1_312 ( .A(_3022__bF_buf3), .B(_3037_), .Y(_1242__6_) );
	INVX1 INVX1_754 ( .A(micro_hash_synth_1_W_0__7_), .Y(_3038_) );
	NOR2X1 NOR2X1_313 ( .A(_3022__bF_buf2), .B(_3038_), .Y(_1242__7_) );
	INVX1 INVX1_755 ( .A(micro_hash_synth_1_W_2__0_), .Y(_3039_) );
	NOR2X1 NOR2X1_314 ( .A(_3022__bF_buf1), .B(_3039_), .Y(_1242__16_) );
	INVX1 INVX1_756 ( .A(micro_hash_synth_1_W_2__1_), .Y(_3040_) );
	NOR2X1 NOR2X1_315 ( .A(_3022__bF_buf0), .B(_3040_), .Y(_1242__17_) );
	INVX1 INVX1_757 ( .A(micro_hash_synth_1_W_2__2_), .Y(_3041_) );
	NOR2X1 NOR2X1_316 ( .A(_3022__bF_buf5), .B(_3041_), .Y(_1242__18_) );
	INVX1 INVX1_758 ( .A(micro_hash_synth_1_W_2__3_), .Y(_3042_) );
	NOR2X1 NOR2X1_317 ( .A(_3022__bF_buf4), .B(_3042_), .Y(_1242__19_) );
	INVX1 INVX1_759 ( .A(micro_hash_synth_1_W_2__4_), .Y(_3043_) );
	NOR2X1 NOR2X1_318 ( .A(_3022__bF_buf3), .B(_3043_), .Y(_1242__20_) );
	INVX1 INVX1_760 ( .A(micro_hash_synth_1_W_2__5_), .Y(_3044_) );
	NOR2X1 NOR2X1_319 ( .A(_3022__bF_buf2), .B(_3044_), .Y(_1242__21_) );
	INVX1 INVX1_761 ( .A(micro_hash_synth_1_W_2__6_), .Y(_3045_) );
	NOR2X1 NOR2X1_320 ( .A(_3022__bF_buf1), .B(_3045_), .Y(_1242__22_) );
	INVX1 INVX1_762 ( .A(micro_hash_synth_1_W_2__7_), .Y(_3046_) );
	NOR2X1 NOR2X1_321 ( .A(_3022__bF_buf0), .B(_3046_), .Y(_1242__23_) );
	NOR2X1 NOR2X1_322 ( .A(_3022__bF_buf5), .B(_3006_), .Y(_1242__24_) );
	NOR2X1 NOR2X1_323 ( .A(_3022__bF_buf4), .B(_3008_), .Y(_1242__25_) );
	NOR2X1 NOR2X1_324 ( .A(_3022__bF_buf3), .B(_3010_), .Y(_1242__26_) );
	NOR2X1 NOR2X1_325 ( .A(_3022__bF_buf2), .B(_3012_), .Y(_1242__27_) );
	NOR2X1 NOR2X1_326 ( .A(_3022__bF_buf1), .B(_3014_), .Y(_1242__28_) );
	NOR2X1 NOR2X1_327 ( .A(_3022__bF_buf0), .B(_3016_), .Y(_1242__29_) );
	NOR2X1 NOR2X1_328 ( .A(_3022__bF_buf5), .B(_3018_), .Y(_1242__30_) );
	NOR2X1 NOR2X1_329 ( .A(_3022__bF_buf4), .B(_3020_), .Y(_1242__31_) );
	INVX1 INVX1_763 ( .A(Hhash_synth1_8_), .Y(_1500_) );
	NOR2X1 NOR2X1_330 ( .A(concatenador_counter_4_), .B(_2927_), .Y(_1501_) );
	INVX1 INVX1_764 ( .A(_1501_), .Y(_1502_) );
	INVX1 INVX1_765 ( .A(concatenador_counter_5_), .Y(_1503_) );
	NOR2X1 NOR2X1_331 ( .A(_1__bF_buf2), .B(_1503_), .Y(_1504_) );
	NAND2X1 NAND2X1_425 ( .A(concatenador_counter_0_bF_buf0), .B(_1504_), .Y(_1505_) );
	NOR2X1 NOR2X1_332 ( .A(_1505_), .B(_1502_), .Y(_1506_) );
	INVX2 INVX2_5 ( .A(_1506__bF_buf3), .Y(_1507_) );
	NOR2X1 NOR2X1_333 ( .A(_3022__bF_buf3), .B(_1507_), .Y(_1508_) );
	NAND3X1 NAND3X1_146 ( .A(reset_L_bF_buf3), .B(_2929_), .C(_1507_), .Y(_1509_) );
	INVX4 INVX4_4 ( .A(_1508_), .Y(_1510_) );
	OAI21X1 OAI21X1_838 ( .A(_1510_), .B(micro_hash_synth_1_b_0_), .C(_1509_), .Y(_1511_) );
	INVX1 INVX1_766 ( .A(micro_hash_synth_1_b_0_), .Y(_1512_) );
	NOR2X1 NOR2X1_334 ( .A(_1500_), .B(_1512_), .Y(_1513_) );
	AOI22X1 AOI22X1_27 ( .A(_1508_), .B(_1513_), .C(_1511_), .D(_1500_), .Y(_1237__8_) );
	INVX1 INVX1_767 ( .A(Hhash_synth1_9_), .Y(_1514_) );
	INVX1 INVX1_768 ( .A(micro_hash_synth_1_b_1_), .Y(_1515_) );
	NOR2X1 NOR2X1_335 ( .A(_1514_), .B(_1515_), .Y(_1516_) );
	NOR2X1 NOR2X1_336 ( .A(Hhash_synth1_9_), .B(micro_hash_synth_1_b_1_), .Y(_1517_) );
	NOR2X1 NOR2X1_337 ( .A(_1517_), .B(_1516_), .Y(_1518_) );
	NAND2X1 NAND2X1_426 ( .A(_1513_), .B(_1518_), .Y(_1519_) );
	OR2X2 OR2X2_39 ( .A(_1518_), .B(_1513_), .Y(_1520_) );
	AOI21X1 AOI21X1_642 ( .A(_1519_), .B(_1520_), .C(_1507_), .Y(_1521_) );
	OAI21X1 OAI21X1_839 ( .A(_2927_), .B(_2921_), .C(reset_L_bF_buf2), .Y(_1522_) );
	INVX4 INVX4_5 ( .A(_1522__bF_buf3), .Y(_1523_) );
	NAND2X1 NAND2X1_427 ( .A(Hhash_synth1_9_), .B(_1523__bF_buf3), .Y(_1524_) );
	AOI21X1 AOI21X1_643 ( .A(_1524_), .B(_1510_), .C(_1521_), .Y(_1237__9_) );
	OAI21X1 OAI21X1_840 ( .A(_1514_), .B(_1515_), .C(_1519_), .Y(_1525_) );
	AND2X2 AND2X2_54 ( .A(Hhash_synth1_10_), .B(micro_hash_synth_1_b_2_), .Y(_1526_) );
	NOR2X1 NOR2X1_338 ( .A(Hhash_synth1_10_), .B(micro_hash_synth_1_b_2_), .Y(_1527_) );
	NOR2X1 NOR2X1_339 ( .A(_1527_), .B(_1526_), .Y(_1528_) );
	XNOR2X1 XNOR2X1_27 ( .A(_1525_), .B(_1528_), .Y(_1529_) );
	NAND2X1 NAND2X1_428 ( .A(Hhash_synth1_10_), .B(_1523__bF_buf2), .Y(_1530_) );
	AOI22X1 AOI22X1_28 ( .A(_1506__bF_buf2), .B(_1529_), .C(_1510_), .D(_1530_), .Y(_1237__10_) );
	AOI21X1 AOI21X1_644 ( .A(_1528_), .B(_1525_), .C(_1526_), .Y(_1531_) );
	INVX1 INVX1_769 ( .A(Hhash_synth1_11_), .Y(_1532_) );
	INVX1 INVX1_770 ( .A(micro_hash_synth_1_b_3_), .Y(_1533_) );
	NOR2X1 NOR2X1_340 ( .A(_1532_), .B(_1533_), .Y(_1534_) );
	NOR2X1 NOR2X1_341 ( .A(Hhash_synth1_11_), .B(micro_hash_synth_1_b_3_), .Y(_1535_) );
	NOR2X1 NOR2X1_342 ( .A(_1535_), .B(_1534_), .Y(_1536_) );
	XOR2X1 XOR2X1_38 ( .A(_1531_), .B(_1536_), .Y(_1537_) );
	OAI21X1 OAI21X1_841 ( .A(Hhash_synth1_11_), .B(_1522__bF_buf2), .C(_1510_), .Y(_1538_) );
	OAI21X1 OAI21X1_842 ( .A(_1507_), .B(_1537_), .C(_1538_), .Y(_1237__11_) );
	XOR2X1 XOR2X1_39 ( .A(Hhash_synth1_12_), .B(micro_hash_synth_1_b_4_), .Y(_1539_) );
	INVX1 INVX1_771 ( .A(_1534_), .Y(_1540_) );
	OAI21X1 OAI21X1_843 ( .A(_1531_), .B(_1535_), .C(_1540_), .Y(_1541_) );
	XNOR2X1 XNOR2X1_28 ( .A(_1541_), .B(_1539_), .Y(_1542_) );
	AOI21X1 AOI21X1_645 ( .A(Hhash_synth1_12_), .B(_1523__bF_buf1), .C(_1508_), .Y(_1543_) );
	AOI21X1 AOI21X1_646 ( .A(_1506__bF_buf1), .B(_1542_), .C(_1543_), .Y(_1237__12_) );
	AOI21X1 AOI21X1_647 ( .A(Hhash_synth1_13_), .B(_1523__bF_buf0), .C(_1508_), .Y(_1544_) );
	AND2X2 AND2X2_55 ( .A(_1541_), .B(_1539_), .Y(_1545_) );
	AOI21X1 AOI21X1_648 ( .A(Hhash_synth1_12_), .B(micro_hash_synth_1_b_4_), .C(_1545_), .Y(_1546_) );
	NAND2X1 NAND2X1_429 ( .A(Hhash_synth1_13_), .B(micro_hash_synth_1_b_5_), .Y(_1547_) );
	INVX1 INVX1_772 ( .A(_1547_), .Y(_1548_) );
	NOR2X1 NOR2X1_343 ( .A(Hhash_synth1_13_), .B(micro_hash_synth_1_b_5_), .Y(_1549_) );
	NOR2X1 NOR2X1_344 ( .A(_1549_), .B(_1548_), .Y(_1550_) );
	XOR2X1 XOR2X1_40 ( .A(_1546_), .B(_1550_), .Y(_1551_) );
	AOI21X1 AOI21X1_649 ( .A(_1506__bF_buf0), .B(_1551_), .C(_1544_), .Y(_1237__13_) );
	XOR2X1 XOR2X1_41 ( .A(Hhash_synth1_14_), .B(micro_hash_synth_1_b_6_), .Y(_1552_) );
	OAI21X1 OAI21X1_844 ( .A(_1546_), .B(_1549_), .C(_1547_), .Y(_1553_) );
	XNOR2X1 XNOR2X1_29 ( .A(_1553_), .B(_1552_), .Y(_1554_) );
	AOI21X1 AOI21X1_650 ( .A(Hhash_synth1_14_), .B(_1523__bF_buf3), .C(_1508_), .Y(_1555_) );
	AOI21X1 AOI21X1_651 ( .A(_1506__bF_buf3), .B(_1554_), .C(_1555_), .Y(_1237__14_) );
	OAI21X1 OAI21X1_845 ( .A(Hhash_synth1_15_), .B(_1522__bF_buf1), .C(_1510_), .Y(_1556_) );
	AND2X2 AND2X2_56 ( .A(Hhash_synth1_14_), .B(micro_hash_synth_1_b_6_), .Y(_1557_) );
	AOI21X1 AOI21X1_652 ( .A(_1552_), .B(_1553_), .C(_1557_), .Y(_1558_) );
	XNOR2X1 XNOR2X1_30 ( .A(Hhash_synth1_15_), .B(micro_hash_synth_1_b_7_), .Y(_1559_) );
	NOR2X1 NOR2X1_345 ( .A(_1559_), .B(_1558_), .Y(_1560_) );
	NAND2X1 NAND2X1_430 ( .A(_1559_), .B(_1558_), .Y(_1561_) );
	NAND2X1 NAND2X1_431 ( .A(_1506__bF_buf2), .B(_1561_), .Y(_1562_) );
	OAI21X1 OAI21X1_846 ( .A(_1562_), .B(_1560_), .C(_1556_), .Y(_1237__15_) );
	INVX1 INVX1_773 ( .A(Hhash_synth1_0_), .Y(_1563_) );
	OAI21X1 OAI21X1_847 ( .A(_1510_), .B(micro_hash_synth_1_a_0_), .C(_1509_), .Y(_1564_) );
	INVX1 INVX1_774 ( .A(micro_hash_synth_1_a_0_), .Y(_1565_) );
	NOR2X1 NOR2X1_346 ( .A(_1563_), .B(_1565_), .Y(_1566_) );
	AOI22X1 AOI22X1_29 ( .A(_1508_), .B(_1566_), .C(_1564_), .D(_1563_), .Y(_1237__0_) );
	INVX1 INVX1_775 ( .A(Hhash_synth1_1_), .Y(_1567_) );
	INVX1 INVX1_776 ( .A(micro_hash_synth_1_a_1_), .Y(_1568_) );
	NOR2X1 NOR2X1_347 ( .A(_1567_), .B(_1568_), .Y(_1569_) );
	NOR2X1 NOR2X1_348 ( .A(Hhash_synth1_1_), .B(micro_hash_synth_1_a_1_), .Y(_1570_) );
	NOR2X1 NOR2X1_349 ( .A(_1570_), .B(_1569_), .Y(_1571_) );
	NAND2X1 NAND2X1_432 ( .A(_1566_), .B(_1571_), .Y(_1572_) );
	OR2X2 OR2X2_40 ( .A(_1571_), .B(_1566_), .Y(_1573_) );
	AOI21X1 AOI21X1_653 ( .A(_1572_), .B(_1573_), .C(_1507_), .Y(_1574_) );
	NAND2X1 NAND2X1_433 ( .A(Hhash_synth1_1_), .B(_1523__bF_buf2), .Y(_1575_) );
	AOI21X1 AOI21X1_654 ( .A(_1575_), .B(_1510_), .C(_1574_), .Y(_1237__1_) );
	OAI21X1 OAI21X1_848 ( .A(_1567_), .B(_1568_), .C(_1572_), .Y(_1576_) );
	AND2X2 AND2X2_57 ( .A(Hhash_synth1_2_), .B(micro_hash_synth_1_a_2_), .Y(_1577_) );
	NOR2X1 NOR2X1_350 ( .A(Hhash_synth1_2_), .B(micro_hash_synth_1_a_2_), .Y(_1578_) );
	NOR2X1 NOR2X1_351 ( .A(_1578_), .B(_1577_), .Y(_1579_) );
	XNOR2X1 XNOR2X1_31 ( .A(_1576_), .B(_1579_), .Y(_1580_) );
	NAND2X1 NAND2X1_434 ( .A(Hhash_synth1_2_), .B(_1523__bF_buf1), .Y(_1581_) );
	AOI22X1 AOI22X1_30 ( .A(_1506__bF_buf1), .B(_1580_), .C(_1510_), .D(_1581_), .Y(_1237__2_) );
	NAND2X1 NAND2X1_435 ( .A(Hhash_synth1_3_), .B(_1523__bF_buf0), .Y(_1582_) );
	AOI21X1 AOI21X1_655 ( .A(_1579_), .B(_1576_), .C(_1577_), .Y(_1583_) );
	AND2X2 AND2X2_58 ( .A(Hhash_synth1_3_), .B(micro_hash_synth_1_a_3_), .Y(_1584_) );
	NOR2X1 NOR2X1_352 ( .A(Hhash_synth1_3_), .B(micro_hash_synth_1_a_3_), .Y(_1585_) );
	NOR2X1 NOR2X1_353 ( .A(_1585_), .B(_1584_), .Y(_1586_) );
	XOR2X1 XOR2X1_42 ( .A(_1583_), .B(_1586_), .Y(_1587_) );
	AOI22X1 AOI22X1_31 ( .A(_1506__bF_buf0), .B(_1587_), .C(_1510_), .D(_1582_), .Y(_1237__3_) );
	XOR2X1 XOR2X1_43 ( .A(Hhash_synth1_4_), .B(micro_hash_synth_1_a_4_), .Y(_1588_) );
	INVX1 INVX1_777 ( .A(_1584_), .Y(_1589_) );
	OAI21X1 OAI21X1_849 ( .A(_1583_), .B(_1585_), .C(_1589_), .Y(_1590_) );
	XNOR2X1 XNOR2X1_32 ( .A(_1590_), .B(_1588_), .Y(_1591_) );
	AOI21X1 AOI21X1_656 ( .A(Hhash_synth1_4_), .B(_1523__bF_buf3), .C(_1508_), .Y(_1592_) );
	AOI21X1 AOI21X1_657 ( .A(_1506__bF_buf3), .B(_1591_), .C(_1592_), .Y(_1237__4_) );
	AOI21X1 AOI21X1_658 ( .A(Hhash_synth1_5_), .B(_1523__bF_buf2), .C(_1508_), .Y(_1593_) );
	AND2X2 AND2X2_59 ( .A(_1590_), .B(_1588_), .Y(_1594_) );
	AOI21X1 AOI21X1_659 ( .A(Hhash_synth1_4_), .B(micro_hash_synth_1_a_4_), .C(_1594_), .Y(_1595_) );
	NAND2X1 NAND2X1_436 ( .A(Hhash_synth1_5_), .B(micro_hash_synth_1_a_5_), .Y(_1596_) );
	INVX1 INVX1_778 ( .A(_1596_), .Y(_1597_) );
	NOR2X1 NOR2X1_354 ( .A(Hhash_synth1_5_), .B(micro_hash_synth_1_a_5_), .Y(_1598_) );
	NOR2X1 NOR2X1_355 ( .A(_1598_), .B(_1597_), .Y(_1599_) );
	OAI21X1 OAI21X1_850 ( .A(_1595_), .B(_1599_), .C(_1506__bF_buf2), .Y(_1600_) );
	AOI21X1 AOI21X1_660 ( .A(_1595_), .B(_1599_), .C(_1600_), .Y(_1601_) );
	NOR2X1 NOR2X1_356 ( .A(_1593_), .B(_1601_), .Y(_1237__5_) );
	XOR2X1 XOR2X1_44 ( .A(Hhash_synth1_6_), .B(micro_hash_synth_1_a_6_), .Y(_1602_) );
	OAI21X1 OAI21X1_851 ( .A(_1595_), .B(_1598_), .C(_1596_), .Y(_1603_) );
	XNOR2X1 XNOR2X1_33 ( .A(_1603_), .B(_1602_), .Y(_1604_) );
	AOI21X1 AOI21X1_661 ( .A(Hhash_synth1_6_), .B(_1523__bF_buf1), .C(_1508_), .Y(_1605_) );
	AOI21X1 AOI21X1_662 ( .A(_1506__bF_buf1), .B(_1604_), .C(_1605_), .Y(_1237__6_) );
	AOI21X1 AOI21X1_663 ( .A(Hhash_synth1_7_), .B(_1523__bF_buf0), .C(_1508_), .Y(_1606_) );
	INVX1 INVX1_779 ( .A(Hhash_synth1_6_), .Y(_1607_) );
	INVX1 INVX1_780 ( .A(micro_hash_synth_1_a_6_), .Y(_1608_) );
	NAND2X1 NAND2X1_437 ( .A(_1602_), .B(_1603_), .Y(_1609_) );
	OAI21X1 OAI21X1_852 ( .A(_1607_), .B(_1608_), .C(_1609_), .Y(_1610_) );
	XNOR2X1 XNOR2X1_34 ( .A(Hhash_synth1_7_), .B(micro_hash_synth_1_a_7_), .Y(_1611_) );
	OAI21X1 OAI21X1_853 ( .A(_1610_), .B(_1611_), .C(_1506__bF_buf0), .Y(_1612_) );
	AOI21X1 AOI21X1_664 ( .A(_1610_), .B(_1611_), .C(_1612_), .Y(_1613_) );
	NOR2X1 NOR2X1_357 ( .A(_1606_), .B(_1613_), .Y(_1237__7_) );
	OAI21X1 OAI21X1_854 ( .A(_2927_), .B(concatenador_counter_4_), .C(concatenador_counter_5_), .Y(_1614_) );
	NOR2X1 NOR2X1_358 ( .A(_3022__bF_buf2), .B(_1614__bF_buf3), .Y(_1615_) );
	INVX4 INVX4_6 ( .A(_1615_), .Y(_1616_) );
	OR2X2 OR2X2_41 ( .A(_1616_), .B(micro_hash_synth_1_k_0_), .Y(_1241__0_) );
	INVX1 INVX1_781 ( .A(micro_hash_synth_1_k_1_), .Y(_1617_) );
	NOR2X1 NOR2X1_359 ( .A(_1617_), .B(_1616_), .Y(_1241__1_) );
	INVX1 INVX1_782 ( .A(micro_hash_synth_1_k_2_), .Y(_1618_) );
	NOR2X1 NOR2X1_360 ( .A(_1618_), .B(_1616_), .Y(_1241__2_) );
	INVX1 INVX1_783 ( .A(micro_hash_synth_1_k_3_), .Y(_1619_) );
	NOR2X1 NOR2X1_361 ( .A(concatenador_counter_0_bF_buf13), .B(concatenador_counter_5_), .Y(_1620_) );
	AOI21X1 AOI21X1_665 ( .A(_1620_), .B(_2926_), .C(_2920_), .Y(_1621_) );
	INVX1 INVX1_784 ( .A(_1621_), .Y(_1622_) );
	NOR2X1 NOR2X1_362 ( .A(_3022__bF_buf1), .B(_1622_), .Y(_1623_) );
	OAI21X1 OAI21X1_855 ( .A(_1614__bF_buf2), .B(_1619_), .C(_1623_), .Y(_1241__3_) );
	INVX1 INVX1_785 ( .A(micro_hash_synth_1_k_4_), .Y(_1624_) );
	OAI21X1 OAI21X1_856 ( .A(_1614__bF_buf1), .B(_1624_), .C(_1623_), .Y(_1241__4_) );
	INVX1 INVX1_786 ( .A(micro_hash_synth_1_k_5_), .Y(_1625_) );
	INVX2 INVX2_6 ( .A(_1614__bF_buf0), .Y(_1626_) );
	INVX2 INVX2_7 ( .A(_1623_), .Y(_1627_) );
	AOI21X1 AOI21X1_666 ( .A(_1625_), .B(_1626_), .C(_1627_), .Y(_1241__5_) );
	AND2X2 AND2X2_60 ( .A(_1615_), .B(micro_hash_synth_1_k_6_), .Y(_1241__6_) );
	OR2X2 OR2X2_42 ( .A(_1616_), .B(micro_hash_synth_1_k_7_), .Y(_1241__7_) );
	INVX1 INVX1_787 ( .A(micro_hash_synth_1_c_0_), .Y(_1628_) );
	INVX4 INVX4_7 ( .A(concatenador_counter_1_bF_buf3), .Y(_1629_) );
	NOR2X1 NOR2X1_363 ( .A(concatenador_counter_2_), .B(_1629__bF_buf3), .Y(_1630_) );
	INVX1 INVX1_788 ( .A(concatenador_counter_2_), .Y(_1631_) );
	NOR2X1 NOR2X1_364 ( .A(concatenador_counter_1_bF_buf2), .B(_1631_), .Y(_1632_) );
	NOR2X1 NOR2X1_365 ( .A(_1630__bF_buf4), .B(_1632__bF_buf4), .Y(_1633_) );
	NOR2X1 NOR2X1_366 ( .A(micro_hash_synth_1_W_5__0_), .B(_2923__bF_buf5), .Y(_1634_) );
	OAI21X1 OAI21X1_857 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_4__0_), .C(concatenador_counter_1_bF_buf1), .Y(_1635_) );
	NOR2X1 NOR2X1_367 ( .A(concatenador_counter_0_bF_buf11), .B(micro_hash_synth_1_W_6__0_), .Y(_1636_) );
	OAI21X1 OAI21X1_858 ( .A(_2923__bF_buf4), .B(micro_hash_synth_1_W_7__0_), .C(_1629__bF_buf2), .Y(_1637_) );
	OAI22X1 OAI22X1_261 ( .A(_1634_), .B(_1635_), .C(_1637_), .D(_1636_), .Y(_1638_) );
	NAND2X1 NAND2X1_438 ( .A(_1633__bF_buf5), .B(_1638_), .Y(_1639_) );
	NAND3X1 NAND3X1_147 ( .A(concatenador_counter_3_), .B(_1629__bF_buf1), .C(_1631_), .Y(_1640_) );
	INVX1 INVX1_789 ( .A(concatenador_counter_3_), .Y(_1641_) );
	OAI21X1 OAI21X1_859 ( .A(concatenador_counter_1_bF_buf0), .B(concatenador_counter_2_), .C(_1641_), .Y(_1642_) );
	NAND2X1 NAND2X1_439 ( .A(_1642_), .B(_1640_), .Y(_1643_) );
	NAND2X1 NAND2X1_440 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_1__0_), .Y(_1644_) );
	OAI21X1 OAI21X1_860 ( .A(_3031_), .B(concatenador_counter_0_bF_buf9), .C(_1644_), .Y(_1645_) );
	NAND2X1 NAND2X1_441 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_3__0_), .Y(_1646_) );
	OAI21X1 OAI21X1_861 ( .A(_3039_), .B(concatenador_counter_0_bF_buf7), .C(_1646_), .Y(_1647_) );
	AOI22X1 AOI22X1_32 ( .A(_1645_), .B(_1630__bF_buf3), .C(_1632__bF_buf3), .D(_1647_), .Y(_1648_) );
	NAND3X1 NAND3X1_148 ( .A(_1643__bF_buf3), .B(_1648_), .C(_1639_), .Y(_1649_) );
	XOR2X1 XOR2X1_45 ( .A(_2926_), .B(concatenador_counter_4_), .Y(_1650_) );
	NOR2X1 NOR2X1_368 ( .A(micro_hash_synth_1_W_13__0_), .B(_2923__bF_buf3), .Y(_1651_) );
	OAI21X1 OAI21X1_862 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_12__0_), .C(concatenador_counter_1_bF_buf7), .Y(_1652_) );
	NOR2X1 NOR2X1_369 ( .A(concatenador_counter_0_bF_buf5), .B(micro_hash_synth_1_W_14__0_), .Y(_1653_) );
	OAI21X1 OAI21X1_863 ( .A(_2923__bF_buf2), .B(micro_hash_synth_1_W_15__0_), .C(_1629__bF_buf0), .Y(_1654_) );
	OAI22X1 OAI22X1_262 ( .A(_1651_), .B(_1652_), .C(_1654_), .D(_1653_), .Y(_1655_) );
	NAND2X1 NAND2X1_442 ( .A(_1633__bF_buf4), .B(_1655_), .Y(_1656_) );
	NAND2X1 NAND2X1_443 ( .A(concatenador_counter_1_bF_buf6), .B(_1631_), .Y(_1657_) );
	NAND2X1 NAND2X1_444 ( .A(concatenador_counter_2_), .B(_1629__bF_buf3), .Y(_1658_) );
	MUX2X1 MUX2X1_15 ( .A(micro_hash_synth_1_W_11__0_), .B(micro_hash_synth_1_W_10__0_), .S(concatenador_counter_0_bF_buf4), .Y(_1659_) );
	MUX2X1 MUX2X1_16 ( .A(micro_hash_synth_1_W_9__0_), .B(micro_hash_synth_1_W_8__0_), .S(concatenador_counter_0_bF_buf3), .Y(_1660_) );
	OAI22X1 OAI22X1_263 ( .A(_1659_), .B(_1658_), .C(_1657_), .D(_1660_), .Y(_1661_) );
	NOR2X1 NOR2X1_370 ( .A(_1643__bF_buf2), .B(_1661_), .Y(_1662_) );
	AOI21X1 AOI21X1_667 ( .A(_1656_), .B(_1662_), .C(_1650_), .Y(_1663_) );
	NOR2X1 NOR2X1_371 ( .A(micro_hash_synth_1_W_21__0_), .B(_2923__bF_buf1), .Y(_1664_) );
	OAI21X1 OAI21X1_864 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_20__0_), .C(concatenador_counter_1_bF_buf5), .Y(_1665_) );
	NOR2X1 NOR2X1_372 ( .A(concatenador_counter_0_bF_buf1), .B(micro_hash_synth_1_W_22__0_), .Y(_1666_) );
	OAI21X1 OAI21X1_865 ( .A(_2923__bF_buf0), .B(micro_hash_synth_1_W_23__0_), .C(_1629__bF_buf2), .Y(_1667_) );
	OAI22X1 OAI22X1_264 ( .A(_1664_), .B(_1665_), .C(_1667_), .D(_1666_), .Y(_1668_) );
	NAND2X1 NAND2X1_445 ( .A(_1633__bF_buf3), .B(_1668_), .Y(_1669_) );
	INVX1 INVX1_790 ( .A(micro_hash_synth_1_W_18__0_), .Y(_1670_) );
	NAND2X1 NAND2X1_446 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_19__0_), .Y(_1671_) );
	OAI21X1 OAI21X1_866 ( .A(_1670_), .B(concatenador_counter_0_bF_buf13), .C(_1671_), .Y(_1672_) );
	INVX1 INVX1_791 ( .A(micro_hash_synth_1_W_16__0_), .Y(_1673_) );
	NAND2X1 NAND2X1_447 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_17__0_), .Y(_1674_) );
	OAI21X1 OAI21X1_867 ( .A(_1673_), .B(concatenador_counter_0_bF_buf11), .C(_1674_), .Y(_1675_) );
	AOI22X1 AOI22X1_33 ( .A(_1672_), .B(_1632__bF_buf2), .C(_1630__bF_buf2), .D(_1675_), .Y(_1676_) );
	NAND3X1 NAND3X1_149 ( .A(_1643__bF_buf1), .B(_1676_), .C(_1669_), .Y(_1677_) );
	OAI21X1 OAI21X1_868 ( .A(concatenador_counter_1_bF_buf4), .B(concatenador_counter_2_), .C(concatenador_counter_3_), .Y(_1678_) );
	OAI21X1 OAI21X1_869 ( .A(_2919_), .B(concatenador_counter_1_bF_buf3), .C(_1678_), .Y(_1679_) );
	XNOR2X1 XNOR2X1_35 ( .A(_2926_), .B(concatenador_counter_4_), .Y(_1680_) );
	MUX2X1 MUX2X1_17 ( .A(micro_hash_synth_1_W_29__0_), .B(micro_hash_synth_1_W_28__0_), .S(concatenador_counter_0_bF_buf10), .Y(_1681_) );
	MUX2X1 MUX2X1_18 ( .A(micro_hash_synth_1_W_31__0_), .B(micro_hash_synth_1_W_30__0_), .S(concatenador_counter_0_bF_buf9), .Y(_1682_) );
	MUX2X1 MUX2X1_19 ( .A(_1682_), .B(_1681_), .S(_1629__bF_buf1), .Y(_1683_) );
	MUX2X1 MUX2X1_20 ( .A(micro_hash_synth_1_W_25__0_), .B(micro_hash_synth_1_W_24__0_), .S(concatenador_counter_0_bF_buf8), .Y(_1684_) );
	MUX2X1 MUX2X1_21 ( .A(micro_hash_synth_1_W_27__0_), .B(micro_hash_synth_1_W_26__0_), .S(concatenador_counter_0_bF_buf7), .Y(_1685_) );
	OAI22X1 OAI22X1_265 ( .A(_1684_), .B(_1657_), .C(_1658_), .D(_1685_), .Y(_1686_) );
	AOI21X1 AOI21X1_668 ( .A(_1633__bF_buf2), .B(_1683_), .C(_1686_), .Y(_1687_) );
	AOI21X1 AOI21X1_669 ( .A(_1679__bF_buf3), .B(_1687_), .C(_1680_), .Y(_1688_) );
	AOI22X1 AOI22X1_34 ( .A(_1663_), .B(_1649_), .C(_1688_), .D(_1677_), .Y(_1689_) );
	INVX1 INVX1_792 ( .A(_1689_), .Y(_1690_) );
	NAND2X1 NAND2X1_448 ( .A(micro_hash_synth_1_k_0_), .B(micro_hash_synth_1_x_0_), .Y(_1691_) );
	INVX1 INVX1_793 ( .A(_1691_), .Y(_1692_) );
	NOR2X1 NOR2X1_373 ( .A(micro_hash_synth_1_k_0_), .B(micro_hash_synth_1_x_0_), .Y(_1693_) );
	NOR2X1 NOR2X1_374 ( .A(_1693_), .B(_1692_), .Y(_1694_) );
	OAI21X1 OAI21X1_870 ( .A(_2927_), .B(_2921_), .C(_1614__bF_buf3), .Y(_1695_) );
	AOI21X1 AOI21X1_670 ( .A(_1694_), .B(_1690_), .C(_1695_), .Y(_1696_) );
	OAI21X1 OAI21X1_871 ( .A(_1690_), .B(_1694_), .C(_1696_), .Y(_1697_) );
	OAI22X1 OAI22X1_266 ( .A(_1628_), .B(_1616_), .C(_1697_), .D(_3022__bF_buf0), .Y(_1240__0_) );
	OAI21X1 OAI21X1_872 ( .A(_1689_), .B(_1693_), .C(_1691_), .Y(_1698_) );
	NOR2X1 NOR2X1_375 ( .A(micro_hash_synth_1_W_21__1_), .B(_2923__bF_buf7), .Y(_1699_) );
	OAI21X1 OAI21X1_873 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_20__1_), .C(concatenador_counter_1_bF_buf2), .Y(_1700_) );
	MUX2X1 MUX2X1_22 ( .A(micro_hash_synth_1_W_23__1_), .B(micro_hash_synth_1_W_22__1_), .S(concatenador_counter_0_bF_buf5), .Y(_1701_) );
	OAI22X1 OAI22X1_267 ( .A(_1701_), .B(concatenador_counter_1_bF_buf1), .C(_1699_), .D(_1700_), .Y(_1702_) );
	INVX1 INVX1_794 ( .A(micro_hash_synth_1_W_18__1_), .Y(_1703_) );
	NAND2X1 NAND2X1_449 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_19__1_), .Y(_1704_) );
	OAI21X1 OAI21X1_874 ( .A(_1703_), .B(concatenador_counter_0_bF_buf3), .C(_1704_), .Y(_1705_) );
	NAND2X1 NAND2X1_450 ( .A(_1632__bF_buf1), .B(_1705_), .Y(_1706_) );
	INVX1 INVX1_795 ( .A(micro_hash_synth_1_W_16__1_), .Y(_1707_) );
	NAND2X1 NAND2X1_451 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_17__1_), .Y(_1708_) );
	OAI21X1 OAI21X1_875 ( .A(_1707_), .B(concatenador_counter_0_bF_buf1), .C(_1708_), .Y(_1709_) );
	NAND2X1 NAND2X1_452 ( .A(_1630__bF_buf1), .B(_1709_), .Y(_1710_) );
	NAND3X1 NAND3X1_150 ( .A(_1643__bF_buf0), .B(_1706_), .C(_1710_), .Y(_1711_) );
	AOI21X1 AOI21X1_671 ( .A(_1633__bF_buf1), .B(_1702_), .C(_1711_), .Y(_1712_) );
	NAND2X1 NAND2X1_453 ( .A(_1657_), .B(_1658_), .Y(_1713_) );
	INVX1 INVX1_796 ( .A(micro_hash_synth_1_W_29__1_), .Y(_1714_) );
	NAND2X1 NAND2X1_454 ( .A(concatenador_counter_0_bF_buf0), .B(_1714_), .Y(_1715_) );
	OR2X2 OR2X2_43 ( .A(concatenador_counter_0_bF_buf13), .B(micro_hash_synth_1_W_28__1_), .Y(_1716_) );
	NAND3X1 NAND3X1_151 ( .A(concatenador_counter_1_bF_buf0), .B(_1716_), .C(_1715_), .Y(_1717_) );
	OR2X2 OR2X2_44 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_30__1_), .Y(_1718_) );
	INVX1 INVX1_797 ( .A(micro_hash_synth_1_W_31__1_), .Y(_1719_) );
	NAND2X1 NAND2X1_455 ( .A(concatenador_counter_0_bF_buf11), .B(_1719_), .Y(_1720_) );
	NAND3X1 NAND3X1_152 ( .A(_1629__bF_buf0), .B(_1718_), .C(_1720_), .Y(_1721_) );
	AOI21X1 AOI21X1_672 ( .A(_1717_), .B(_1721_), .C(_1713_), .Y(_1722_) );
	INVX1 INVX1_798 ( .A(micro_hash_synth_1_W_24__1_), .Y(_1723_) );
	NAND2X1 NAND2X1_456 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_25__1_), .Y(_1724_) );
	OAI21X1 OAI21X1_876 ( .A(_1723_), .B(concatenador_counter_0_bF_buf9), .C(_1724_), .Y(_1725_) );
	NAND2X1 NAND2X1_457 ( .A(_1630__bF_buf0), .B(_1725_), .Y(_1726_) );
	NAND2X1 NAND2X1_458 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_27__1_), .Y(_1727_) );
	OAI21X1 OAI21X1_877 ( .A(_2933_), .B(concatenador_counter_0_bF_buf7), .C(_1727_), .Y(_1728_) );
	NAND2X1 NAND2X1_459 ( .A(_1632__bF_buf0), .B(_1728_), .Y(_1729_) );
	NAND3X1 NAND3X1_153 ( .A(_1679__bF_buf2), .B(_1726_), .C(_1729_), .Y(_1730_) );
	OAI21X1 OAI21X1_878 ( .A(_1730_), .B(_1722_), .C(_1650_), .Y(_1731_) );
	NOR2X1 NOR2X1_376 ( .A(micro_hash_synth_1_W_13__1_), .B(_2923__bF_buf6), .Y(_1732_) );
	OAI21X1 OAI21X1_879 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_12__1_), .C(concatenador_counter_1_bF_buf7), .Y(_1733_) );
	MUX2X1 MUX2X1_23 ( .A(micro_hash_synth_1_W_15__1_), .B(micro_hash_synth_1_W_14__1_), .S(concatenador_counter_0_bF_buf5), .Y(_1734_) );
	OAI22X1 OAI22X1_268 ( .A(_1734_), .B(concatenador_counter_1_bF_buf6), .C(_1732_), .D(_1733_), .Y(_1735_) );
	INVX1 INVX1_799 ( .A(micro_hash_synth_1_W_10__1_), .Y(_1736_) );
	NAND2X1 NAND2X1_460 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_11__1_), .Y(_1737_) );
	OAI21X1 OAI21X1_880 ( .A(_1736_), .B(concatenador_counter_0_bF_buf3), .C(_1737_), .Y(_1738_) );
	NAND2X1 NAND2X1_461 ( .A(_1632__bF_buf4), .B(_1738_), .Y(_1739_) );
	NAND2X1 NAND2X1_462 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_9__1_), .Y(_1740_) );
	OAI21X1 OAI21X1_881 ( .A(_2992_), .B(concatenador_counter_0_bF_buf1), .C(_1740_), .Y(_1741_) );
	NAND2X1 NAND2X1_463 ( .A(_1630__bF_buf4), .B(_1741_), .Y(_1742_) );
	NAND3X1 NAND3X1_154 ( .A(_1679__bF_buf1), .B(_1739_), .C(_1742_), .Y(_1743_) );
	AOI21X1 AOI21X1_673 ( .A(_1633__bF_buf0), .B(_1735_), .C(_1743_), .Y(_1744_) );
	INVX1 INVX1_800 ( .A(micro_hash_synth_1_W_5__1_), .Y(_1745_) );
	NAND2X1 NAND2X1_464 ( .A(concatenador_counter_0_bF_buf0), .B(_1745_), .Y(_1746_) );
	OR2X2 OR2X2_45 ( .A(concatenador_counter_0_bF_buf13), .B(micro_hash_synth_1_W_4__1_), .Y(_1747_) );
	NAND3X1 NAND3X1_155 ( .A(concatenador_counter_1_bF_buf5), .B(_1747_), .C(_1746_), .Y(_1748_) );
	OR2X2 OR2X2_46 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_6__1_), .Y(_1749_) );
	INVX1 INVX1_801 ( .A(micro_hash_synth_1_W_7__1_), .Y(_1750_) );
	NAND2X1 NAND2X1_465 ( .A(concatenador_counter_0_bF_buf11), .B(_1750_), .Y(_1751_) );
	NAND3X1 NAND3X1_156 ( .A(_1629__bF_buf3), .B(_1749_), .C(_1751_), .Y(_1752_) );
	AOI21X1 AOI21X1_674 ( .A(_1748_), .B(_1752_), .C(_1713_), .Y(_1753_) );
	NAND2X1 NAND2X1_466 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_1__1_), .Y(_1754_) );
	OAI21X1 OAI21X1_882 ( .A(_3032_), .B(concatenador_counter_0_bF_buf9), .C(_1754_), .Y(_1755_) );
	NAND2X1 NAND2X1_467 ( .A(_1630__bF_buf3), .B(_1755_), .Y(_1756_) );
	NAND2X1 NAND2X1_468 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_3__1_), .Y(_1757_) );
	OAI21X1 OAI21X1_883 ( .A(_3040_), .B(concatenador_counter_0_bF_buf7), .C(_1757_), .Y(_1758_) );
	NAND2X1 NAND2X1_469 ( .A(_1632__bF_buf3), .B(_1758_), .Y(_1759_) );
	NAND3X1 NAND3X1_157 ( .A(_1643__bF_buf3), .B(_1756_), .C(_1759_), .Y(_1760_) );
	OAI21X1 OAI21X1_884 ( .A(_1760_), .B(_1753_), .C(_1680_), .Y(_1761_) );
	OAI22X1 OAI22X1_269 ( .A(_1731_), .B(_1712_), .C(_1744_), .D(_1761_), .Y(_1762_) );
	AND2X2 AND2X2_61 ( .A(micro_hash_synth_1_k_1_), .B(micro_hash_synth_1_x_1_), .Y(_1763_) );
	NOR2X1 NOR2X1_377 ( .A(micro_hash_synth_1_k_1_), .B(micro_hash_synth_1_x_1_), .Y(_1764_) );
	NOR2X1 NOR2X1_378 ( .A(_1764_), .B(_1763_), .Y(_1765_) );
	NAND2X1 NAND2X1_470 ( .A(_1765_), .B(_1762_), .Y(_1766_) );
	NAND2X1 NAND2X1_471 ( .A(_1633__bF_buf5), .B(_1702_), .Y(_1767_) );
	AOI21X1 AOI21X1_675 ( .A(_1630__bF_buf2), .B(_1709_), .C(_1679__bF_buf0), .Y(_1768_) );
	NAND3X1 NAND3X1_158 ( .A(_1706_), .B(_1768_), .C(_1767_), .Y(_1769_) );
	NOR2X1 NOR2X1_379 ( .A(micro_hash_synth_1_W_29__1_), .B(_2923__bF_buf5), .Y(_1770_) );
	OAI21X1 OAI21X1_885 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_28__1_), .C(concatenador_counter_1_bF_buf4), .Y(_1771_) );
	MUX2X1 MUX2X1_24 ( .A(micro_hash_synth_1_W_31__1_), .B(micro_hash_synth_1_W_30__1_), .S(concatenador_counter_0_bF_buf5), .Y(_1772_) );
	OAI22X1 OAI22X1_270 ( .A(_1772_), .B(concatenador_counter_1_bF_buf3), .C(_1770_), .D(_1771_), .Y(_1773_) );
	NAND2X1 NAND2X1_472 ( .A(_1633__bF_buf4), .B(_1773_), .Y(_1774_) );
	AOI21X1 AOI21X1_676 ( .A(_1632__bF_buf2), .B(_1728_), .C(_1643__bF_buf2), .Y(_1775_) );
	NAND3X1 NAND3X1_159 ( .A(_1726_), .B(_1775_), .C(_1774_), .Y(_1776_) );
	NAND3X1 NAND3X1_160 ( .A(_1650_), .B(_1769_), .C(_1776_), .Y(_1777_) );
	NAND2X1 NAND2X1_473 ( .A(_1633__bF_buf3), .B(_1735_), .Y(_1778_) );
	AOI21X1 AOI21X1_677 ( .A(_1630__bF_buf1), .B(_1741_), .C(_1643__bF_buf1), .Y(_1779_) );
	NAND3X1 NAND3X1_161 ( .A(_1739_), .B(_1779_), .C(_1778_), .Y(_1780_) );
	NOR2X1 NOR2X1_380 ( .A(micro_hash_synth_1_W_5__1_), .B(_2923__bF_buf4), .Y(_1781_) );
	OAI21X1 OAI21X1_886 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_4__1_), .C(concatenador_counter_1_bF_buf2), .Y(_1782_) );
	MUX2X1 MUX2X1_25 ( .A(micro_hash_synth_1_W_7__1_), .B(micro_hash_synth_1_W_6__1_), .S(concatenador_counter_0_bF_buf3), .Y(_1783_) );
	OAI22X1 OAI22X1_271 ( .A(_1783_), .B(concatenador_counter_1_bF_buf1), .C(_1781_), .D(_1782_), .Y(_1784_) );
	NAND2X1 NAND2X1_474 ( .A(_1633__bF_buf2), .B(_1784_), .Y(_1785_) );
	AOI21X1 AOI21X1_678 ( .A(_1632__bF_buf1), .B(_1758_), .C(_1679__bF_buf3), .Y(_1786_) );
	NAND3X1 NAND3X1_162 ( .A(_1756_), .B(_1786_), .C(_1785_), .Y(_1787_) );
	NAND3X1 NAND3X1_163 ( .A(_1680_), .B(_1780_), .C(_1787_), .Y(_1788_) );
	INVX1 INVX1_802 ( .A(_1765_), .Y(_1789_) );
	NAND3X1 NAND3X1_164 ( .A(_1789_), .B(_1777_), .C(_1788_), .Y(_1790_) );
	NAND3X1 NAND3X1_165 ( .A(_1766_), .B(_1790_), .C(_1698_), .Y(_1791_) );
	INVX1 INVX1_803 ( .A(_1791_), .Y(_1792_) );
	INVX2 INVX2_8 ( .A(_1695_), .Y(_1793_) );
	NAND2X1 NAND2X1_475 ( .A(_1790_), .B(_1766_), .Y(_1794_) );
	INVX1 INVX1_804 ( .A(_1794_), .Y(_1795_) );
	OAI21X1 OAI21X1_887 ( .A(_1795_), .B(_1698_), .C(_1793_), .Y(_1796_) );
	AOI21X1 AOI21X1_679 ( .A(micro_hash_synth_1_c_1_), .B(_1626_), .C(_1522__bF_buf0), .Y(_1797_) );
	OAI21X1 OAI21X1_888 ( .A(_1796_), .B(_1792_), .C(_1797_), .Y(_1240__1_) );
	AOI21X1 AOI21X1_680 ( .A(_1777_), .B(_1788_), .C(_1789_), .Y(_1798_) );
	NOR2X1 NOR2X1_381 ( .A(micro_hash_synth_1_W_21__2_), .B(_2923__bF_buf3), .Y(_1799_) );
	OAI21X1 OAI21X1_889 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_20__2_), .C(concatenador_counter_1_bF_buf0), .Y(_1800_) );
	MUX2X1 MUX2X1_26 ( .A(micro_hash_synth_1_W_23__2_), .B(micro_hash_synth_1_W_22__2_), .S(concatenador_counter_0_bF_buf1), .Y(_1801_) );
	OAI22X1 OAI22X1_272 ( .A(_1801_), .B(concatenador_counter_1_bF_buf7), .C(_1799_), .D(_1800_), .Y(_1802_) );
	NAND2X1 NAND2X1_476 ( .A(_1633__bF_buf1), .B(_1802_), .Y(_1803_) );
	INVX1 INVX1_805 ( .A(micro_hash_synth_1_W_18__2_), .Y(_1804_) );
	NAND2X1 NAND2X1_477 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_19__2_), .Y(_1805_) );
	OAI21X1 OAI21X1_890 ( .A(_1804_), .B(concatenador_counter_0_bF_buf13), .C(_1805_), .Y(_1806_) );
	NAND2X1 NAND2X1_478 ( .A(_1632__bF_buf0), .B(_1806_), .Y(_1807_) );
	INVX1 INVX1_806 ( .A(micro_hash_synth_1_W_16__2_), .Y(_1808_) );
	NAND2X1 NAND2X1_479 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_17__2_), .Y(_1809_) );
	OAI21X1 OAI21X1_891 ( .A(_1808_), .B(concatenador_counter_0_bF_buf11), .C(_1809_), .Y(_1810_) );
	AOI21X1 AOI21X1_681 ( .A(_1630__bF_buf0), .B(_1810_), .C(_1679__bF_buf2), .Y(_1811_) );
	NAND3X1 NAND3X1_166 ( .A(_1807_), .B(_1811_), .C(_1803_), .Y(_1812_) );
	NOR2X1 NOR2X1_382 ( .A(micro_hash_synth_1_W_29__2_), .B(_2923__bF_buf2), .Y(_1813_) );
	OAI21X1 OAI21X1_892 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_28__2_), .C(concatenador_counter_1_bF_buf6), .Y(_1814_) );
	NOR2X1 NOR2X1_383 ( .A(concatenador_counter_0_bF_buf9), .B(micro_hash_synth_1_W_30__2_), .Y(_1815_) );
	OAI21X1 OAI21X1_893 ( .A(_2923__bF_buf1), .B(micro_hash_synth_1_W_31__2_), .C(_1629__bF_buf2), .Y(_1816_) );
	OAI22X1 OAI22X1_273 ( .A(_1813_), .B(_1814_), .C(_1816_), .D(_1815_), .Y(_1817_) );
	NAND2X1 NAND2X1_480 ( .A(_1633__bF_buf0), .B(_1817_), .Y(_1818_) );
	INVX1 INVX1_807 ( .A(micro_hash_synth_1_W_24__2_), .Y(_1819_) );
	NAND2X1 NAND2X1_481 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_25__2_), .Y(_1820_) );
	OAI21X1 OAI21X1_894 ( .A(_1819_), .B(concatenador_counter_0_bF_buf7), .C(_1820_), .Y(_1821_) );
	NAND2X1 NAND2X1_482 ( .A(_1630__bF_buf4), .B(_1821_), .Y(_1822_) );
	NAND2X1 NAND2X1_483 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_27__2_), .Y(_1823_) );
	OAI21X1 OAI21X1_895 ( .A(_2938_), .B(concatenador_counter_0_bF_buf5), .C(_1823_), .Y(_1824_) );
	AOI21X1 AOI21X1_682 ( .A(_1632__bF_buf4), .B(_1824_), .C(_1643__bF_buf0), .Y(_1825_) );
	NAND3X1 NAND3X1_167 ( .A(_1822_), .B(_1825_), .C(_1818_), .Y(_1826_) );
	NAND3X1 NAND3X1_168 ( .A(_1650_), .B(_1812_), .C(_1826_), .Y(_1827_) );
	NOR2X1 NOR2X1_384 ( .A(micro_hash_synth_1_W_13__2_), .B(_2923__bF_buf0), .Y(_1828_) );
	OAI21X1 OAI21X1_896 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_12__2_), .C(concatenador_counter_1_bF_buf5), .Y(_1829_) );
	MUX2X1 MUX2X1_27 ( .A(micro_hash_synth_1_W_15__2_), .B(micro_hash_synth_1_W_14__2_), .S(concatenador_counter_0_bF_buf3), .Y(_1830_) );
	OAI22X1 OAI22X1_274 ( .A(_1830_), .B(concatenador_counter_1_bF_buf4), .C(_1828_), .D(_1829_), .Y(_1831_) );
	NAND2X1 NAND2X1_484 ( .A(_1633__bF_buf5), .B(_1831_), .Y(_1832_) );
	NAND2X1 NAND2X1_485 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_9__2_), .Y(_1833_) );
	OAI21X1 OAI21X1_897 ( .A(_2994_), .B(concatenador_counter_0_bF_buf1), .C(_1833_), .Y(_1834_) );
	NAND2X1 NAND2X1_486 ( .A(_1630__bF_buf3), .B(_1834_), .Y(_1835_) );
	INVX1 INVX1_808 ( .A(micro_hash_synth_1_W_10__2_), .Y(_1836_) );
	NAND2X1 NAND2X1_487 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_11__2_), .Y(_1837_) );
	OAI21X1 OAI21X1_898 ( .A(_1836_), .B(concatenador_counter_0_bF_buf13), .C(_1837_), .Y(_1838_) );
	AOI21X1 AOI21X1_683 ( .A(_1632__bF_buf3), .B(_1838_), .C(_1643__bF_buf3), .Y(_1839_) );
	NAND3X1 NAND3X1_169 ( .A(_1835_), .B(_1839_), .C(_1832_), .Y(_1840_) );
	NOR2X1 NOR2X1_385 ( .A(micro_hash_synth_1_W_5__2_), .B(_2923__bF_buf7), .Y(_1841_) );
	OAI21X1 OAI21X1_899 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_4__2_), .C(concatenador_counter_1_bF_buf3), .Y(_1842_) );
	NOR2X1 NOR2X1_386 ( .A(concatenador_counter_0_bF_buf11), .B(micro_hash_synth_1_W_6__2_), .Y(_1843_) );
	OAI21X1 OAI21X1_900 ( .A(_2923__bF_buf6), .B(micro_hash_synth_1_W_7__2_), .C(_1629__bF_buf1), .Y(_1844_) );
	OAI22X1 OAI22X1_275 ( .A(_1841_), .B(_1842_), .C(_1844_), .D(_1843_), .Y(_1845_) );
	NAND2X1 NAND2X1_488 ( .A(_1633__bF_buf4), .B(_1845_), .Y(_1846_) );
	NAND2X1 NAND2X1_489 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_1__2_), .Y(_1847_) );
	OAI21X1 OAI21X1_901 ( .A(_3033_), .B(concatenador_counter_0_bF_buf9), .C(_1847_), .Y(_1848_) );
	NAND2X1 NAND2X1_490 ( .A(_1630__bF_buf2), .B(_1848_), .Y(_1849_) );
	NAND2X1 NAND2X1_491 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_3__2_), .Y(_1850_) );
	OAI21X1 OAI21X1_902 ( .A(_3041_), .B(concatenador_counter_0_bF_buf7), .C(_1850_), .Y(_1851_) );
	AOI21X1 AOI21X1_684 ( .A(_1632__bF_buf2), .B(_1851_), .C(_1679__bF_buf1), .Y(_1852_) );
	NAND3X1 NAND3X1_170 ( .A(_1849_), .B(_1852_), .C(_1846_), .Y(_1853_) );
	NAND3X1 NAND3X1_171 ( .A(_1680_), .B(_1840_), .C(_1853_), .Y(_1854_) );
	NAND2X1 NAND2X1_492 ( .A(micro_hash_synth_1_k_2_), .B(micro_hash_synth_1_x_2_), .Y(_1855_) );
	INVX1 INVX1_809 ( .A(micro_hash_synth_1_x_2_), .Y(_1856_) );
	NAND2X1 NAND2X1_493 ( .A(_1618_), .B(_1856_), .Y(_1857_) );
	AND2X2 AND2X2_62 ( .A(_1857_), .B(_1855_), .Y(_1858_) );
	INVX1 INVX1_810 ( .A(_1858_), .Y(_1859_) );
	AOI21X1 AOI21X1_685 ( .A(_1827_), .B(_1854_), .C(_1859_), .Y(_1860_) );
	NAND2X1 NAND2X1_494 ( .A(_1630__bF_buf1), .B(_1810_), .Y(_1861_) );
	NAND3X1 NAND3X1_172 ( .A(_1643__bF_buf2), .B(_1807_), .C(_1861_), .Y(_1862_) );
	AOI21X1 AOI21X1_686 ( .A(_1633__bF_buf3), .B(_1802_), .C(_1862_), .Y(_1863_) );
	INVX1 INVX1_811 ( .A(micro_hash_synth_1_W_29__2_), .Y(_1864_) );
	NAND2X1 NAND2X1_495 ( .A(concatenador_counter_0_bF_buf6), .B(_1864_), .Y(_1865_) );
	OR2X2 OR2X2_47 ( .A(concatenador_counter_0_bF_buf5), .B(micro_hash_synth_1_W_28__2_), .Y(_1866_) );
	NAND3X1 NAND3X1_173 ( .A(concatenador_counter_1_bF_buf2), .B(_1866_), .C(_1865_), .Y(_1867_) );
	OR2X2 OR2X2_48 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_30__2_), .Y(_1868_) );
	INVX1 INVX1_812 ( .A(micro_hash_synth_1_W_31__2_), .Y(_1869_) );
	NAND2X1 NAND2X1_496 ( .A(concatenador_counter_0_bF_buf3), .B(_1869_), .Y(_1870_) );
	NAND3X1 NAND3X1_174 ( .A(_1629__bF_buf0), .B(_1868_), .C(_1870_), .Y(_1871_) );
	AOI21X1 AOI21X1_687 ( .A(_1867_), .B(_1871_), .C(_1713_), .Y(_1872_) );
	NAND2X1 NAND2X1_497 ( .A(_1632__bF_buf1), .B(_1824_), .Y(_1873_) );
	NAND3X1 NAND3X1_175 ( .A(_1679__bF_buf0), .B(_1822_), .C(_1873_), .Y(_1874_) );
	OAI21X1 OAI21X1_903 ( .A(_1874_), .B(_1872_), .C(_1650_), .Y(_1875_) );
	NAND2X1 NAND2X1_498 ( .A(_1632__bF_buf0), .B(_1838_), .Y(_1876_) );
	NAND3X1 NAND3X1_176 ( .A(_1679__bF_buf3), .B(_1835_), .C(_1876_), .Y(_1877_) );
	AOI21X1 AOI21X1_688 ( .A(_1633__bF_buf2), .B(_1831_), .C(_1877_), .Y(_1878_) );
	INVX1 INVX1_813 ( .A(micro_hash_synth_1_W_5__2_), .Y(_1879_) );
	NAND2X1 NAND2X1_499 ( .A(concatenador_counter_0_bF_buf2), .B(_1879_), .Y(_1880_) );
	OR2X2 OR2X2_49 ( .A(concatenador_counter_0_bF_buf1), .B(micro_hash_synth_1_W_4__2_), .Y(_1881_) );
	NAND3X1 NAND3X1_177 ( .A(concatenador_counter_1_bF_buf1), .B(_1881_), .C(_1880_), .Y(_1882_) );
	OR2X2 OR2X2_50 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_6__2_), .Y(_1883_) );
	INVX1 INVX1_814 ( .A(micro_hash_synth_1_W_7__2_), .Y(_1884_) );
	NAND2X1 NAND2X1_500 ( .A(concatenador_counter_0_bF_buf13), .B(_1884_), .Y(_1885_) );
	NAND3X1 NAND3X1_178 ( .A(_1629__bF_buf3), .B(_1883_), .C(_1885_), .Y(_1886_) );
	AOI21X1 AOI21X1_689 ( .A(_1882_), .B(_1886_), .C(_1713_), .Y(_1887_) );
	NAND2X1 NAND2X1_501 ( .A(_1632__bF_buf4), .B(_1851_), .Y(_1888_) );
	NAND3X1 NAND3X1_179 ( .A(_1643__bF_buf1), .B(_1849_), .C(_1888_), .Y(_1889_) );
	OAI21X1 OAI21X1_904 ( .A(_1889_), .B(_1887_), .C(_1680_), .Y(_1890_) );
	OAI22X1 OAI22X1_276 ( .A(_1875_), .B(_1863_), .C(_1878_), .D(_1890_), .Y(_1891_) );
	NOR2X1 NOR2X1_387 ( .A(_1858_), .B(_1891_), .Y(_1892_) );
	OAI22X1 OAI22X1_277 ( .A(_1763_), .B(_1798_), .C(_1892_), .D(_1860_), .Y(_1893_) );
	AOI21X1 AOI21X1_690 ( .A(_1765_), .B(_1762_), .C(_1763_), .Y(_1894_) );
	NAND2X1 NAND2X1_502 ( .A(_1858_), .B(_1891_), .Y(_1895_) );
	NAND3X1 NAND3X1_180 ( .A(_1859_), .B(_1827_), .C(_1854_), .Y(_1896_) );
	NAND3X1 NAND3X1_181 ( .A(_1895_), .B(_1896_), .C(_1894_), .Y(_1897_) );
	NAND2X1 NAND2X1_503 ( .A(_1893_), .B(_1897_), .Y(_1898_) );
	NOR2X1 NOR2X1_388 ( .A(_1792_), .B(_1898_), .Y(_1899_) );
	AOI21X1 AOI21X1_691 ( .A(_1893_), .B(_1897_), .C(_1791_), .Y(_1900_) );
	INVX1 INVX1_815 ( .A(_1900_), .Y(_1901_) );
	NAND2X1 NAND2X1_504 ( .A(_1793_), .B(_1901_), .Y(_1902_) );
	AOI21X1 AOI21X1_692 ( .A(micro_hash_synth_1_c_2_), .B(_1626_), .C(_1522__bF_buf3), .Y(_1903_) );
	OAI21X1 OAI21X1_905 ( .A(_1902_), .B(_1899_), .C(_1903_), .Y(_1240__2_) );
	NAND2X1 NAND2X1_505 ( .A(_1895_), .B(_1896_), .Y(_1904_) );
	NOR2X1 NOR2X1_389 ( .A(_1894_), .B(_1904_), .Y(_1905_) );
	NOR2X1 NOR2X1_390 ( .A(_1905_), .B(_1900_), .Y(_1906_) );
	AOI21X1 AOI21X1_693 ( .A(micro_hash_synth_1_k_2_), .B(micro_hash_synth_1_x_2_), .C(_1860_), .Y(_1907_) );
	NAND2X1 NAND2X1_506 ( .A(micro_hash_synth_1_k_3_), .B(micro_hash_synth_1_x_3_), .Y(_1908_) );
	INVX1 INVX1_816 ( .A(micro_hash_synth_1_x_3_), .Y(_1909_) );
	NAND2X1 NAND2X1_507 ( .A(_1619_), .B(_1909_), .Y(_1910_) );
	AND2X2 AND2X2_63 ( .A(_1910_), .B(_1908_), .Y(_1911_) );
	INVX1 INVX1_817 ( .A(_1911_), .Y(_1912_) );
	NOR2X1 NOR2X1_391 ( .A(micro_hash_synth_1_W_29__3_), .B(_2923__bF_buf5), .Y(_1913_) );
	OAI21X1 OAI21X1_906 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_28__3_), .C(concatenador_counter_1_bF_buf0), .Y(_1914_) );
	NOR2X1 NOR2X1_392 ( .A(concatenador_counter_0_bF_buf11), .B(micro_hash_synth_1_W_30__3_), .Y(_1915_) );
	OAI21X1 OAI21X1_907 ( .A(_2923__bF_buf4), .B(micro_hash_synth_1_W_31__3_), .C(_1629__bF_buf2), .Y(_1916_) );
	OAI22X1 OAI22X1_278 ( .A(_1913_), .B(_1914_), .C(_1916_), .D(_1915_), .Y(_1917_) );
	NAND2X1 NAND2X1_508 ( .A(_1633__bF_buf1), .B(_1917_), .Y(_1918_) );
	INVX1 INVX1_818 ( .A(micro_hash_synth_1_W_24__3_), .Y(_1919_) );
	NAND2X1 NAND2X1_509 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_25__3_), .Y(_1920_) );
	OAI21X1 OAI21X1_908 ( .A(_1919_), .B(concatenador_counter_0_bF_buf9), .C(_1920_), .Y(_1921_) );
	NAND2X1 NAND2X1_510 ( .A(_1630__bF_buf0), .B(_1921_), .Y(_1922_) );
	NAND2X1 NAND2X1_511 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_27__3_), .Y(_1923_) );
	OAI21X1 OAI21X1_909 ( .A(_2943_), .B(concatenador_counter_0_bF_buf7), .C(_1923_), .Y(_1924_) );
	NAND2X1 NAND2X1_512 ( .A(_1632__bF_buf3), .B(_1924_), .Y(_1925_) );
	AND2X2 AND2X2_64 ( .A(_1922_), .B(_1925_), .Y(_1926_) );
	AOI21X1 AOI21X1_694 ( .A(_1918_), .B(_1926_), .C(_1643__bF_buf0), .Y(_1927_) );
	NOR2X1 NOR2X1_393 ( .A(micro_hash_synth_1_W_21__3_), .B(_2923__bF_buf3), .Y(_1928_) );
	OAI21X1 OAI21X1_910 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_20__3_), .C(concatenador_counter_1_bF_buf7), .Y(_1929_) );
	NOR2X1 NOR2X1_394 ( .A(concatenador_counter_0_bF_buf5), .B(micro_hash_synth_1_W_22__3_), .Y(_1930_) );
	OAI21X1 OAI21X1_911 ( .A(_2923__bF_buf2), .B(micro_hash_synth_1_W_23__3_), .C(_1629__bF_buf1), .Y(_1931_) );
	OAI22X1 OAI22X1_279 ( .A(_1928_), .B(_1929_), .C(_1931_), .D(_1930_), .Y(_1932_) );
	NAND2X1 NAND2X1_513 ( .A(_1633__bF_buf0), .B(_1932_), .Y(_1933_) );
	INVX1 INVX1_819 ( .A(micro_hash_synth_1_W_18__3_), .Y(_1934_) );
	NAND2X1 NAND2X1_514 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_19__3_), .Y(_1935_) );
	OAI21X1 OAI21X1_912 ( .A(_1934_), .B(concatenador_counter_0_bF_buf3), .C(_1935_), .Y(_1936_) );
	NAND2X1 NAND2X1_515 ( .A(_1632__bF_buf2), .B(_1936_), .Y(_1937_) );
	INVX1 INVX1_820 ( .A(micro_hash_synth_1_W_16__3_), .Y(_1938_) );
	NAND2X1 NAND2X1_516 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_17__3_), .Y(_1939_) );
	OAI21X1 OAI21X1_913 ( .A(_1938_), .B(concatenador_counter_0_bF_buf1), .C(_1939_), .Y(_1940_) );
	NAND2X1 NAND2X1_517 ( .A(_1630__bF_buf4), .B(_1940_), .Y(_1941_) );
	AND2X2 AND2X2_65 ( .A(_1937_), .B(_1941_), .Y(_1942_) );
	AOI21X1 AOI21X1_695 ( .A(_1933_), .B(_1942_), .C(_1679__bF_buf2), .Y(_1943_) );
	OAI21X1 OAI21X1_914 ( .A(_1927_), .B(_1943_), .C(_1650_), .Y(_1944_) );
	NOR2X1 NOR2X1_395 ( .A(micro_hash_synth_1_W_13__3_), .B(_2923__bF_buf1), .Y(_1945_) );
	OAI21X1 OAI21X1_915 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_12__3_), .C(concatenador_counter_1_bF_buf6), .Y(_1946_) );
	NOR2X1 NOR2X1_396 ( .A(concatenador_counter_0_bF_buf13), .B(micro_hash_synth_1_W_14__3_), .Y(_1947_) );
	OAI21X1 OAI21X1_916 ( .A(_2923__bF_buf0), .B(micro_hash_synth_1_W_15__3_), .C(_1629__bF_buf0), .Y(_1948_) );
	OAI22X1 OAI22X1_280 ( .A(_1945_), .B(_1946_), .C(_1948_), .D(_1947_), .Y(_1949_) );
	NAND2X1 NAND2X1_518 ( .A(_1633__bF_buf5), .B(_1949_), .Y(_1950_) );
	INVX1 INVX1_821 ( .A(micro_hash_synth_1_W_10__3_), .Y(_1951_) );
	NAND2X1 NAND2X1_519 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_11__3_), .Y(_1952_) );
	OAI21X1 OAI21X1_917 ( .A(_1951_), .B(concatenador_counter_0_bF_buf11), .C(_1952_), .Y(_1953_) );
	NAND2X1 NAND2X1_520 ( .A(_1632__bF_buf1), .B(_1953_), .Y(_1954_) );
	NAND2X1 NAND2X1_521 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_9__3_), .Y(_1955_) );
	OAI21X1 OAI21X1_918 ( .A(_2996_), .B(concatenador_counter_0_bF_buf9), .C(_1955_), .Y(_1956_) );
	AOI21X1 AOI21X1_696 ( .A(_1630__bF_buf3), .B(_1956_), .C(_1643__bF_buf3), .Y(_1957_) );
	NAND3X1 NAND3X1_182 ( .A(_1954_), .B(_1957_), .C(_1950_), .Y(_1958_) );
	NOR2X1 NOR2X1_397 ( .A(micro_hash_synth_1_W_5__3_), .B(_2923__bF_buf7), .Y(_1959_) );
	OAI21X1 OAI21X1_919 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_4__3_), .C(concatenador_counter_1_bF_buf5), .Y(_1960_) );
	MUX2X1 MUX2X1_28 ( .A(micro_hash_synth_1_W_7__3_), .B(micro_hash_synth_1_W_6__3_), .S(concatenador_counter_0_bF_buf7), .Y(_1961_) );
	OAI22X1 OAI22X1_281 ( .A(_1961_), .B(concatenador_counter_1_bF_buf4), .C(_1959_), .D(_1960_), .Y(_1962_) );
	AND2X2 AND2X2_66 ( .A(_1962_), .B(_1633__bF_buf4), .Y(_1963_) );
	NAND2X1 NAND2X1_522 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_1__3_), .Y(_1964_) );
	OAI21X1 OAI21X1_920 ( .A(_3034_), .B(concatenador_counter_0_bF_buf5), .C(_1964_), .Y(_1965_) );
	NAND2X1 NAND2X1_523 ( .A(_1630__bF_buf2), .B(_1965_), .Y(_1966_) );
	NAND2X1 NAND2X1_524 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_3__3_), .Y(_1967_) );
	OAI21X1 OAI21X1_921 ( .A(_3042_), .B(concatenador_counter_0_bF_buf3), .C(_1967_), .Y(_1968_) );
	NAND2X1 NAND2X1_525 ( .A(_1632__bF_buf0), .B(_1968_), .Y(_1969_) );
	NAND3X1 NAND3X1_183 ( .A(_1643__bF_buf2), .B(_1966_), .C(_1969_), .Y(_1970_) );
	OR2X2 OR2X2_51 ( .A(_1963_), .B(_1970_), .Y(_1971_) );
	NAND3X1 NAND3X1_184 ( .A(_1680_), .B(_1958_), .C(_1971_), .Y(_1972_) );
	NAND3X1 NAND3X1_185 ( .A(_1912_), .B(_1944_), .C(_1972_), .Y(_1973_) );
	AND2X2 AND2X2_67 ( .A(_1932_), .B(_1633__bF_buf3), .Y(_1974_) );
	NAND3X1 NAND3X1_186 ( .A(_1643__bF_buf1), .B(_1937_), .C(_1941_), .Y(_1975_) );
	AND2X2 AND2X2_68 ( .A(_1917_), .B(_1633__bF_buf2), .Y(_1976_) );
	NAND3X1 NAND3X1_187 ( .A(_1679__bF_buf1), .B(_1922_), .C(_1925_), .Y(_1977_) );
	OAI22X1 OAI22X1_282 ( .A(_1974_), .B(_1975_), .C(_1976_), .D(_1977_), .Y(_1978_) );
	NAND2X1 NAND2X1_526 ( .A(_1650_), .B(_1978_), .Y(_1979_) );
	AND2X2 AND2X2_69 ( .A(_1949_), .B(_1633__bF_buf1), .Y(_1980_) );
	NAND2X1 NAND2X1_527 ( .A(_1630__bF_buf1), .B(_1956_), .Y(_1981_) );
	NAND3X1 NAND3X1_188 ( .A(_1679__bF_buf0), .B(_1954_), .C(_1981_), .Y(_1982_) );
	OAI22X1 OAI22X1_283 ( .A(_1963_), .B(_1970_), .C(_1980_), .D(_1982_), .Y(_1983_) );
	NAND2X1 NAND2X1_528 ( .A(_1680_), .B(_1983_), .Y(_1984_) );
	NAND3X1 NAND3X1_189 ( .A(_1911_), .B(_1984_), .C(_1979_), .Y(_1985_) );
	NAND2X1 NAND2X1_529 ( .A(_1985_), .B(_1973_), .Y(_1986_) );
	NAND2X1 NAND2X1_530 ( .A(_1907_), .B(_1986_), .Y(_1987_) );
	OR2X2 OR2X2_52 ( .A(_1986_), .B(_1907_), .Y(_1988_) );
	NAND2X1 NAND2X1_531 ( .A(_1987_), .B(_1988_), .Y(_1989_) );
	AOI21X1 AOI21X1_697 ( .A(_1989_), .B(_1906_), .C(_1695_), .Y(_1990_) );
	OAI21X1 OAI21X1_922 ( .A(_1906_), .B(_1989_), .C(_1990_), .Y(_1991_) );
	AOI21X1 AOI21X1_698 ( .A(micro_hash_synth_1_c_3_), .B(_1626_), .C(_1522__bF_buf2), .Y(_1992_) );
	NAND2X1 NAND2X1_532 ( .A(_1992_), .B(_1991_), .Y(_1240__3_) );
	AND2X2 AND2X2_70 ( .A(_1985_), .B(_1908_), .Y(_1993_) );
	INVX1 INVX1_822 ( .A(micro_hash_synth_1_x_4_), .Y(_1994_) );
	NOR2X1 NOR2X1_398 ( .A(_1624_), .B(_1994_), .Y(_1995_) );
	NOR2X1 NOR2X1_399 ( .A(micro_hash_synth_1_k_4_), .B(micro_hash_synth_1_x_4_), .Y(_1996_) );
	NOR2X1 NOR2X1_400 ( .A(_1996_), .B(_1995_), .Y(_1997_) );
	NOR2X1 NOR2X1_401 ( .A(micro_hash_synth_1_W_29__4_), .B(_2923__bF_buf6), .Y(_1998_) );
	OAI21X1 OAI21X1_923 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_28__4_), .C(concatenador_counter_1_bF_buf3), .Y(_1999_) );
	NOR2X1 NOR2X1_402 ( .A(concatenador_counter_0_bF_buf1), .B(micro_hash_synth_1_W_30__4_), .Y(_2000_) );
	OAI21X1 OAI21X1_924 ( .A(_2923__bF_buf5), .B(micro_hash_synth_1_W_31__4_), .C(_1629__bF_buf3), .Y(_2001_) );
	OAI22X1 OAI22X1_284 ( .A(_1998_), .B(_1999_), .C(_2001_), .D(_2000_), .Y(_2002_) );
	INVX1 INVX1_823 ( .A(micro_hash_synth_1_W_24__4_), .Y(_2003_) );
	NAND2X1 NAND2X1_533 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_25__4_), .Y(_2004_) );
	OAI21X1 OAI21X1_925 ( .A(_2003_), .B(concatenador_counter_0_bF_buf13), .C(_2004_), .Y(_2005_) );
	NAND2X1 NAND2X1_534 ( .A(_1630__bF_buf0), .B(_2005_), .Y(_2006_) );
	NAND2X1 NAND2X1_535 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_27__4_), .Y(_2007_) );
	OAI21X1 OAI21X1_926 ( .A(_2946_), .B(concatenador_counter_0_bF_buf11), .C(_2007_), .Y(_2008_) );
	NAND2X1 NAND2X1_536 ( .A(_1632__bF_buf4), .B(_2008_), .Y(_2009_) );
	NAND3X1 NAND3X1_190 ( .A(_1679__bF_buf3), .B(_2006_), .C(_2009_), .Y(_2010_) );
	AOI21X1 AOI21X1_699 ( .A(_1633__bF_buf0), .B(_2002_), .C(_2010_), .Y(_2011_) );
	NOR2X1 NOR2X1_403 ( .A(micro_hash_synth_1_W_13__4_), .B(_2923__bF_buf4), .Y(_2012_) );
	OAI21X1 OAI21X1_927 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_12__4_), .C(concatenador_counter_1_bF_buf2), .Y(_2013_) );
	NOR2X1 NOR2X1_404 ( .A(concatenador_counter_0_bF_buf9), .B(micro_hash_synth_1_W_14__4_), .Y(_2014_) );
	OAI21X1 OAI21X1_928 ( .A(_2923__bF_buf3), .B(micro_hash_synth_1_W_15__4_), .C(_1629__bF_buf2), .Y(_2015_) );
	OAI22X1 OAI22X1_285 ( .A(_2012_), .B(_2013_), .C(_2015_), .D(_2014_), .Y(_2016_) );
	INVX1 INVX1_824 ( .A(micro_hash_synth_1_W_10__4_), .Y(_2017_) );
	NAND2X1 NAND2X1_537 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_11__4_), .Y(_2018_) );
	OAI21X1 OAI21X1_929 ( .A(_2017_), .B(concatenador_counter_0_bF_buf7), .C(_2018_), .Y(_2019_) );
	NAND2X1 NAND2X1_538 ( .A(_1632__bF_buf3), .B(_2019_), .Y(_2020_) );
	NAND2X1 NAND2X1_539 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_9__4_), .Y(_2021_) );
	OAI21X1 OAI21X1_930 ( .A(_2998_), .B(concatenador_counter_0_bF_buf5), .C(_2021_), .Y(_2022_) );
	NAND2X1 NAND2X1_540 ( .A(_1630__bF_buf4), .B(_2022_), .Y(_2023_) );
	NAND3X1 NAND3X1_191 ( .A(_1679__bF_buf2), .B(_2020_), .C(_2023_), .Y(_2024_) );
	AOI21X1 AOI21X1_700 ( .A(_1633__bF_buf5), .B(_2016_), .C(_2024_), .Y(_2025_) );
	NOR2X1 NOR2X1_405 ( .A(micro_hash_synth_1_W_21__4_), .B(_2923__bF_buf2), .Y(_2026_) );
	OAI21X1 OAI21X1_931 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_20__4_), .C(concatenador_counter_1_bF_buf1), .Y(_2027_) );
	MUX2X1 MUX2X1_29 ( .A(micro_hash_synth_1_W_23__4_), .B(micro_hash_synth_1_W_22__4_), .S(concatenador_counter_0_bF_buf3), .Y(_2028_) );
	OAI22X1 OAI22X1_286 ( .A(_2028_), .B(concatenador_counter_1_bF_buf0), .C(_2026_), .D(_2027_), .Y(_2029_) );
	AND2X2 AND2X2_71 ( .A(_2029_), .B(_1633__bF_buf4), .Y(_2030_) );
	INVX1 INVX1_825 ( .A(micro_hash_synth_1_W_18__4_), .Y(_2031_) );
	NAND2X1 NAND2X1_541 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_19__4_), .Y(_2032_) );
	OAI21X1 OAI21X1_932 ( .A(_2031_), .B(concatenador_counter_0_bF_buf1), .C(_2032_), .Y(_2033_) );
	NAND2X1 NAND2X1_542 ( .A(_1632__bF_buf2), .B(_2033_), .Y(_2034_) );
	INVX1 INVX1_826 ( .A(micro_hash_synth_1_W_16__4_), .Y(_2035_) );
	NAND2X1 NAND2X1_543 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_17__4_), .Y(_2036_) );
	OAI21X1 OAI21X1_933 ( .A(_2035_), .B(concatenador_counter_0_bF_buf13), .C(_2036_), .Y(_2037_) );
	NAND2X1 NAND2X1_544 ( .A(_1630__bF_buf3), .B(_2037_), .Y(_2038_) );
	NAND3X1 NAND3X1_192 ( .A(_1643__bF_buf0), .B(_2034_), .C(_2038_), .Y(_2039_) );
	OAI21X1 OAI21X1_934 ( .A(_2030_), .B(_2039_), .C(_1650_), .Y(_2040_) );
	NOR2X1 NOR2X1_406 ( .A(micro_hash_synth_1_W_5__4_), .B(_2923__bF_buf1), .Y(_2041_) );
	OAI21X1 OAI21X1_935 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_4__4_), .C(concatenador_counter_1_bF_buf7), .Y(_2042_) );
	MUX2X1 MUX2X1_30 ( .A(micro_hash_synth_1_W_7__4_), .B(micro_hash_synth_1_W_6__4_), .S(concatenador_counter_0_bF_buf11), .Y(_2043_) );
	OAI22X1 OAI22X1_287 ( .A(_2043_), .B(concatenador_counter_1_bF_buf6), .C(_2041_), .D(_2042_), .Y(_2044_) );
	AND2X2 AND2X2_72 ( .A(_2044_), .B(_1633__bF_buf3), .Y(_2045_) );
	NAND2X1 NAND2X1_545 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_1__4_), .Y(_2046_) );
	OAI21X1 OAI21X1_936 ( .A(_3035_), .B(concatenador_counter_0_bF_buf9), .C(_2046_), .Y(_2047_) );
	NAND2X1 NAND2X1_546 ( .A(_1630__bF_buf2), .B(_2047_), .Y(_2048_) );
	NAND2X1 NAND2X1_547 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_3__4_), .Y(_2049_) );
	OAI21X1 OAI21X1_937 ( .A(_3043_), .B(concatenador_counter_0_bF_buf7), .C(_2049_), .Y(_2050_) );
	NAND2X1 NAND2X1_548 ( .A(_1632__bF_buf1), .B(_2050_), .Y(_2051_) );
	NAND3X1 NAND3X1_193 ( .A(_1643__bF_buf3), .B(_2048_), .C(_2051_), .Y(_2052_) );
	OAI21X1 OAI21X1_938 ( .A(_2045_), .B(_2052_), .C(_1680_), .Y(_2053_) );
	OAI22X1 OAI22X1_288 ( .A(_2040_), .B(_2011_), .C(_2025_), .D(_2053_), .Y(_2054_) );
	NOR2X1 NOR2X1_407 ( .A(_1997_), .B(_2054_), .Y(_2055_) );
	INVX1 INVX1_827 ( .A(_1997_), .Y(_2056_) );
	NAND2X1 NAND2X1_549 ( .A(_1633__bF_buf2), .B(_2002_), .Y(_2057_) );
	AND2X2 AND2X2_73 ( .A(_2006_), .B(_2009_), .Y(_2058_) );
	AOI21X1 AOI21X1_701 ( .A(_2057_), .B(_2058_), .C(_1643__bF_buf2), .Y(_2059_) );
	NAND2X1 NAND2X1_550 ( .A(_1633__bF_buf1), .B(_2029_), .Y(_2060_) );
	AND2X2 AND2X2_74 ( .A(_2034_), .B(_2038_), .Y(_2061_) );
	AOI21X1 AOI21X1_702 ( .A(_2060_), .B(_2061_), .C(_1679__bF_buf1), .Y(_2062_) );
	OAI21X1 OAI21X1_939 ( .A(_2059_), .B(_2062_), .C(_1650_), .Y(_2063_) );
	NAND2X1 NAND2X1_551 ( .A(_1633__bF_buf0), .B(_2016_), .Y(_2064_) );
	AND2X2 AND2X2_75 ( .A(_2020_), .B(_2023_), .Y(_2065_) );
	AOI21X1 AOI21X1_703 ( .A(_2064_), .B(_2065_), .C(_1643__bF_buf1), .Y(_2066_) );
	NAND2X1 NAND2X1_552 ( .A(_1633__bF_buf5), .B(_2044_), .Y(_2067_) );
	AND2X2 AND2X2_76 ( .A(_2048_), .B(_2051_), .Y(_2068_) );
	AOI21X1 AOI21X1_704 ( .A(_2067_), .B(_2068_), .C(_1679__bF_buf0), .Y(_2069_) );
	OAI21X1 OAI21X1_940 ( .A(_2066_), .B(_2069_), .C(_1680_), .Y(_2070_) );
	AOI21X1 AOI21X1_705 ( .A(_2063_), .B(_2070_), .C(_2056_), .Y(_2071_) );
	OAI21X1 OAI21X1_941 ( .A(_2055_), .B(_2071_), .C(_1993_), .Y(_2072_) );
	OAI21X1 OAI21X1_942 ( .A(_1619_), .B(_1909_), .C(_1985_), .Y(_2073_) );
	NOR2X1 NOR2X1_408 ( .A(_2071_), .B(_2055_), .Y(_2074_) );
	NAND2X1 NAND2X1_553 ( .A(_2073_), .B(_2074_), .Y(_2075_) );
	NAND2X1 NAND2X1_554 ( .A(_2075_), .B(_2072_), .Y(_2076_) );
	OAI22X1 OAI22X1_289 ( .A(_1894_), .B(_1904_), .C(_1986_), .D(_1907_), .Y(_2077_) );
	OAI21X1 OAI21X1_943 ( .A(_1900_), .B(_2077_), .C(_1987_), .Y(_2078_) );
	AND2X2 AND2X2_77 ( .A(_2078_), .B(_2076_), .Y(_2079_) );
	OAI21X1 OAI21X1_944 ( .A(_2078_), .B(_2076_), .C(_1793_), .Y(_2080_) );
	AOI21X1 AOI21X1_706 ( .A(micro_hash_synth_1_c_4_), .B(_1626_), .C(_1522__bF_buf1), .Y(_2081_) );
	OAI21X1 OAI21X1_945 ( .A(_2079_), .B(_2080_), .C(_2081_), .Y(_1240__4_) );
	OAI21X1 OAI21X1_946 ( .A(_2078_), .B(_2076_), .C(_2075_), .Y(_2082_) );
	XOR2X1 XOR2X1_46 ( .A(micro_hash_synth_1_k_5_), .B(micro_hash_synth_1_x_5_), .Y(_2083_) );
	MUX2X1 MUX2X1_31 ( .A(micro_hash_synth_1_W_21__5_), .B(micro_hash_synth_1_W_20__5_), .S(concatenador_counter_0_bF_buf6), .Y(_2084_) );
	MUX2X1 MUX2X1_32 ( .A(micro_hash_synth_1_W_23__5_), .B(micro_hash_synth_1_W_22__5_), .S(concatenador_counter_0_bF_buf5), .Y(_2085_) );
	MUX2X1 MUX2X1_33 ( .A(_2085_), .B(_2084_), .S(_1629__bF_buf1), .Y(_2086_) );
	AND2X2 AND2X2_78 ( .A(_2086_), .B(_1633__bF_buf4), .Y(_2087_) );
	INVX1 INVX1_828 ( .A(micro_hash_synth_1_W_18__5_), .Y(_2088_) );
	NAND2X1 NAND2X1_555 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_19__5_), .Y(_2089_) );
	OAI21X1 OAI21X1_947 ( .A(_2088_), .B(concatenador_counter_0_bF_buf3), .C(_2089_), .Y(_2090_) );
	NAND2X1 NAND2X1_556 ( .A(_1632__bF_buf0), .B(_2090_), .Y(_2091_) );
	INVX1 INVX1_829 ( .A(micro_hash_synth_1_W_16__5_), .Y(_2092_) );
	NAND2X1 NAND2X1_557 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_17__5_), .Y(_2093_) );
	OAI21X1 OAI21X1_948 ( .A(_2092_), .B(concatenador_counter_0_bF_buf1), .C(_2093_), .Y(_2094_) );
	NAND2X1 NAND2X1_558 ( .A(_1630__bF_buf1), .B(_2094_), .Y(_2095_) );
	NAND3X1 NAND3X1_194 ( .A(_1643__bF_buf0), .B(_2091_), .C(_2095_), .Y(_2096_) );
	NOR2X1 NOR2X1_409 ( .A(micro_hash_synth_1_W_29__5_), .B(_2923__bF_buf0), .Y(_2097_) );
	OAI21X1 OAI21X1_949 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_28__5_), .C(concatenador_counter_1_bF_buf5), .Y(_2098_) );
	MUX2X1 MUX2X1_34 ( .A(micro_hash_synth_1_W_31__5_), .B(micro_hash_synth_1_W_30__5_), .S(concatenador_counter_0_bF_buf13), .Y(_2099_) );
	OAI22X1 OAI22X1_290 ( .A(_2099_), .B(concatenador_counter_1_bF_buf4), .C(_2097_), .D(_2098_), .Y(_2100_) );
	AND2X2 AND2X2_79 ( .A(_2100_), .B(_1633__bF_buf3), .Y(_2101_) );
	NAND2X1 NAND2X1_559 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_27__5_), .Y(_2102_) );
	OAI21X1 OAI21X1_950 ( .A(_2949_), .B(concatenador_counter_0_bF_buf11), .C(_2102_), .Y(_2103_) );
	NAND2X1 NAND2X1_560 ( .A(_1632__bF_buf4), .B(_2103_), .Y(_2104_) );
	INVX1 INVX1_830 ( .A(micro_hash_synth_1_W_24__5_), .Y(_2105_) );
	NAND2X1 NAND2X1_561 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_25__5_), .Y(_2106_) );
	OAI21X1 OAI21X1_951 ( .A(_2105_), .B(concatenador_counter_0_bF_buf9), .C(_2106_), .Y(_2107_) );
	NAND2X1 NAND2X1_562 ( .A(_1630__bF_buf0), .B(_2107_), .Y(_2108_) );
	NAND3X1 NAND3X1_195 ( .A(_1679__bF_buf3), .B(_2104_), .C(_2108_), .Y(_2109_) );
	OAI22X1 OAI22X1_291 ( .A(_2087_), .B(_2096_), .C(_2101_), .D(_2109_), .Y(_2110_) );
	NAND2X1 NAND2X1_563 ( .A(_1650_), .B(_2110_), .Y(_2111_) );
	MUX2X1 MUX2X1_35 ( .A(micro_hash_synth_1_W_13__5_), .B(micro_hash_synth_1_W_12__5_), .S(concatenador_counter_0_bF_buf8), .Y(_2112_) );
	MUX2X1 MUX2X1_36 ( .A(micro_hash_synth_1_W_15__5_), .B(micro_hash_synth_1_W_14__5_), .S(concatenador_counter_0_bF_buf7), .Y(_2113_) );
	MUX2X1 MUX2X1_37 ( .A(_2113_), .B(_2112_), .S(_1629__bF_buf0), .Y(_2114_) );
	AND2X2 AND2X2_80 ( .A(_2114_), .B(_1633__bF_buf2), .Y(_2115_) );
	NAND2X1 NAND2X1_564 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_9__5_), .Y(_2116_) );
	OAI21X1 OAI21X1_952 ( .A(_3000_), .B(concatenador_counter_0_bF_buf5), .C(_2116_), .Y(_2117_) );
	NAND2X1 NAND2X1_565 ( .A(_1630__bF_buf4), .B(_2117_), .Y(_2118_) );
	INVX1 INVX1_831 ( .A(micro_hash_synth_1_W_10__5_), .Y(_2119_) );
	NAND2X1 NAND2X1_566 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_11__5_), .Y(_2120_) );
	OAI21X1 OAI21X1_953 ( .A(_2119_), .B(concatenador_counter_0_bF_buf3), .C(_2120_), .Y(_2121_) );
	NAND2X1 NAND2X1_567 ( .A(_1632__bF_buf3), .B(_2121_), .Y(_2122_) );
	NAND3X1 NAND3X1_196 ( .A(_1679__bF_buf2), .B(_2118_), .C(_2122_), .Y(_2123_) );
	NOR2X1 NOR2X1_410 ( .A(micro_hash_synth_1_W_5__5_), .B(_2923__bF_buf7), .Y(_2124_) );
	OAI21X1 OAI21X1_954 ( .A(concatenador_counter_0_bF_buf2), .B(micro_hash_synth_1_W_4__5_), .C(concatenador_counter_1_bF_buf3), .Y(_2125_) );
	MUX2X1 MUX2X1_38 ( .A(micro_hash_synth_1_W_7__5_), .B(micro_hash_synth_1_W_6__5_), .S(concatenador_counter_0_bF_buf1), .Y(_2126_) );
	OAI22X1 OAI22X1_292 ( .A(_2126_), .B(concatenador_counter_1_bF_buf2), .C(_2124_), .D(_2125_), .Y(_2127_) );
	AND2X2 AND2X2_81 ( .A(_2127_), .B(_1633__bF_buf1), .Y(_2128_) );
	NAND2X1 NAND2X1_568 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_3__5_), .Y(_2129_) );
	OAI21X1 OAI21X1_955 ( .A(_3044_), .B(concatenador_counter_0_bF_buf13), .C(_2129_), .Y(_2130_) );
	NAND2X1 NAND2X1_569 ( .A(_1632__bF_buf2), .B(_2130_), .Y(_2131_) );
	NAND2X1 NAND2X1_570 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_1__5_), .Y(_2132_) );
	OAI21X1 OAI21X1_956 ( .A(_3036_), .B(concatenador_counter_0_bF_buf11), .C(_2132_), .Y(_2133_) );
	NAND2X1 NAND2X1_571 ( .A(_1630__bF_buf3), .B(_2133_), .Y(_2134_) );
	NAND3X1 NAND3X1_197 ( .A(_1643__bF_buf3), .B(_2131_), .C(_2134_), .Y(_2135_) );
	OAI22X1 OAI22X1_293 ( .A(_2115_), .B(_2123_), .C(_2128_), .D(_2135_), .Y(_2136_) );
	NAND2X1 NAND2X1_572 ( .A(_1680_), .B(_2136_), .Y(_2137_) );
	AOI21X1 AOI21X1_707 ( .A(_2111_), .B(_2137_), .C(_2083_), .Y(_2138_) );
	INVX1 INVX1_832 ( .A(_2083_), .Y(_2139_) );
	OR2X2 OR2X2_53 ( .A(_2087_), .B(_2096_), .Y(_2140_) );
	OR2X2 OR2X2_54 ( .A(_2101_), .B(_2109_), .Y(_2141_) );
	NAND3X1 NAND3X1_198 ( .A(_1650_), .B(_2140_), .C(_2141_), .Y(_2142_) );
	OR2X2 OR2X2_55 ( .A(_2115_), .B(_2123_), .Y(_2143_) );
	OR2X2 OR2X2_56 ( .A(_2128_), .B(_2135_), .Y(_2144_) );
	NAND3X1 NAND3X1_199 ( .A(_1680_), .B(_2143_), .C(_2144_), .Y(_2145_) );
	AOI21X1 AOI21X1_708 ( .A(_2142_), .B(_2145_), .C(_2139_), .Y(_2146_) );
	OAI22X1 OAI22X1_294 ( .A(_1995_), .B(_2071_), .C(_2146_), .D(_2138_), .Y(_2147_) );
	AOI21X1 AOI21X1_709 ( .A(_1997_), .B(_2054_), .C(_1995_), .Y(_2148_) );
	NAND3X1 NAND3X1_200 ( .A(_2139_), .B(_2142_), .C(_2145_), .Y(_2149_) );
	NAND3X1 NAND3X1_201 ( .A(_2083_), .B(_2111_), .C(_2137_), .Y(_2150_) );
	NAND3X1 NAND3X1_202 ( .A(_2149_), .B(_2150_), .C(_2148_), .Y(_2151_) );
	NAND2X1 NAND2X1_573 ( .A(_2151_), .B(_2147_), .Y(_2152_) );
	XNOR2X1 XNOR2X1_36 ( .A(_2082_), .B(_2152_), .Y(_2153_) );
	AOI21X1 AOI21X1_710 ( .A(micro_hash_synth_1_c_5_), .B(_1626_), .C(_1522__bF_buf0), .Y(_2154_) );
	OAI21X1 OAI21X1_957 ( .A(_2153_), .B(_1695_), .C(_2154_), .Y(_1240__5_) );
	NAND3X1 NAND3X1_203 ( .A(_2072_), .B(_2075_), .C(_2152_), .Y(_2155_) );
	AND2X2 AND2X2_82 ( .A(_2074_), .B(_2073_), .Y(_2156_) );
	NAND2X1 NAND2X1_574 ( .A(_2150_), .B(_2149_), .Y(_2157_) );
	NOR2X1 NOR2X1_411 ( .A(_2148_), .B(_2157_), .Y(_2158_) );
	AOI21X1 AOI21X1_711 ( .A(_2152_), .B(_2156_), .C(_2158_), .Y(_2159_) );
	OAI21X1 OAI21X1_958 ( .A(_2078_), .B(_2155_), .C(_2159_), .Y(_2160_) );
	AOI21X1 AOI21X1_712 ( .A(micro_hash_synth_1_k_5_), .B(micro_hash_synth_1_x_5_), .C(_2146_), .Y(_2161_) );
	INVX1 INVX1_833 ( .A(_2161_), .Y(_2162_) );
	AND2X2 AND2X2_83 ( .A(micro_hash_synth_1_k_6_), .B(micro_hash_synth_1_x_6_), .Y(_2163_) );
	NOR2X1 NOR2X1_412 ( .A(micro_hash_synth_1_k_6_), .B(micro_hash_synth_1_x_6_), .Y(_2164_) );
	NOR2X1 NOR2X1_413 ( .A(_2164_), .B(_2163_), .Y(_2165_) );
	INVX1 INVX1_834 ( .A(_2165_), .Y(_2166_) );
	NOR2X1 NOR2X1_414 ( .A(micro_hash_synth_1_W_21__6_), .B(_2923__bF_buf6), .Y(_2167_) );
	OAI21X1 OAI21X1_959 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_20__6_), .C(concatenador_counter_1_bF_buf1), .Y(_2168_) );
	AOI21X1 AOI21X1_713 ( .A(concatenador_counter_0_bF_buf9), .B(_2954_), .C(concatenador_counter_1_bF_buf0), .Y(_2169_) );
	OAI21X1 OAI21X1_960 ( .A(concatenador_counter_0_bF_buf8), .B(micro_hash_synth_1_W_22__6_), .C(_2169_), .Y(_2170_) );
	OAI21X1 OAI21X1_961 ( .A(_2167_), .B(_2168_), .C(_2170_), .Y(_2171_) );
	INVX1 INVX1_835 ( .A(micro_hash_synth_1_W_18__6_), .Y(_2172_) );
	AOI21X1 AOI21X1_714 ( .A(_2923__bF_buf5), .B(_2172_), .C(_1658_), .Y(_2173_) );
	OAI21X1 OAI21X1_962 ( .A(_2923__bF_buf4), .B(micro_hash_synth_1_W_19__6_), .C(_2173_), .Y(_2174_) );
	INVX1 INVX1_836 ( .A(micro_hash_synth_1_W_16__6_), .Y(_2175_) );
	AOI21X1 AOI21X1_715 ( .A(_2923__bF_buf3), .B(_2175_), .C(_1657_), .Y(_2176_) );
	OAI21X1 OAI21X1_963 ( .A(_2923__bF_buf2), .B(micro_hash_synth_1_W_17__6_), .C(_2176_), .Y(_2177_) );
	NAND2X1 NAND2X1_575 ( .A(_2174_), .B(_2177_), .Y(_2178_) );
	AOI21X1 AOI21X1_716 ( .A(_1633__bF_buf0), .B(_2171_), .C(_2178_), .Y(_2179_) );
	NOR2X1 NOR2X1_415 ( .A(micro_hash_synth_1_W_29__6_), .B(_2923__bF_buf1), .Y(_2180_) );
	OAI21X1 OAI21X1_964 ( .A(concatenador_counter_0_bF_buf7), .B(micro_hash_synth_1_W_28__6_), .C(concatenador_counter_1_bF_buf7), .Y(_2181_) );
	NOR2X1 NOR2X1_416 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_30__6_), .Y(_2182_) );
	OAI21X1 OAI21X1_965 ( .A(_2923__bF_buf0), .B(micro_hash_synth_1_W_31__6_), .C(_1629__bF_buf3), .Y(_2183_) );
	OAI22X1 OAI22X1_295 ( .A(_2180_), .B(_2181_), .C(_2183_), .D(_2182_), .Y(_2184_) );
	AND2X2 AND2X2_84 ( .A(_2184_), .B(_1633__bF_buf5), .Y(_2185_) );
	INVX1 INVX1_837 ( .A(micro_hash_synth_1_W_24__6_), .Y(_2186_) );
	AOI21X1 AOI21X1_717 ( .A(_2923__bF_buf7), .B(_2186_), .C(_1657_), .Y(_2187_) );
	OAI21X1 OAI21X1_966 ( .A(_2923__bF_buf6), .B(micro_hash_synth_1_W_25__6_), .C(_2187_), .Y(_2188_) );
	AOI21X1 AOI21X1_718 ( .A(_2923__bF_buf5), .B(_2952_), .C(_1658_), .Y(_2189_) );
	OAI21X1 OAI21X1_967 ( .A(_2923__bF_buf4), .B(micro_hash_synth_1_W_27__6_), .C(_2189_), .Y(_2190_) );
	NAND2X1 NAND2X1_576 ( .A(_2188_), .B(_2190_), .Y(_2191_) );
	OAI21X1 OAI21X1_968 ( .A(_2191_), .B(_2185_), .C(_1679__bF_buf1), .Y(_2192_) );
	OAI21X1 OAI21X1_969 ( .A(_1679__bF_buf0), .B(_2179_), .C(_2192_), .Y(_2193_) );
	NAND2X1 NAND2X1_577 ( .A(_1650_), .B(_2193_), .Y(_2194_) );
	NOR2X1 NOR2X1_417 ( .A(micro_hash_synth_1_W_13__6_), .B(_2923__bF_buf3), .Y(_2195_) );
	OAI21X1 OAI21X1_970 ( .A(concatenador_counter_0_bF_buf5), .B(micro_hash_synth_1_W_12__6_), .C(concatenador_counter_1_bF_buf6), .Y(_2196_) );
	INVX1 INVX1_838 ( .A(micro_hash_synth_1_W_15__6_), .Y(_2197_) );
	AOI21X1 AOI21X1_719 ( .A(concatenador_counter_0_bF_buf4), .B(_2197_), .C(concatenador_counter_1_bF_buf5), .Y(_2198_) );
	OAI21X1 OAI21X1_971 ( .A(concatenador_counter_0_bF_buf3), .B(micro_hash_synth_1_W_14__6_), .C(_2198_), .Y(_2199_) );
	OAI21X1 OAI21X1_972 ( .A(_2195_), .B(_2196_), .C(_2199_), .Y(_2200_) );
	AND2X2 AND2X2_85 ( .A(_2200_), .B(_1633__bF_buf4), .Y(_2201_) );
	INVX1 INVX1_839 ( .A(micro_hash_synth_1_W_9__6_), .Y(_2202_) );
	AOI21X1 AOI21X1_720 ( .A(concatenador_counter_0_bF_buf2), .B(_2202_), .C(_1657_), .Y(_2203_) );
	OAI21X1 OAI21X1_973 ( .A(concatenador_counter_0_bF_buf1), .B(micro_hash_synth_1_W_8__6_), .C(_2203_), .Y(_2204_) );
	INVX1 INVX1_840 ( .A(micro_hash_synth_1_W_10__6_), .Y(_2205_) );
	AOI21X1 AOI21X1_721 ( .A(_2923__bF_buf2), .B(_2205_), .C(_1658_), .Y(_2206_) );
	OAI21X1 OAI21X1_974 ( .A(_2923__bF_buf1), .B(micro_hash_synth_1_W_11__6_), .C(_2206_), .Y(_2207_) );
	NAND2X1 NAND2X1_578 ( .A(_2204_), .B(_2207_), .Y(_2208_) );
	OAI21X1 OAI21X1_975 ( .A(_2201_), .B(_2208_), .C(_1679__bF_buf3), .Y(_2209_) );
	NOR2X1 NOR2X1_418 ( .A(micro_hash_synth_1_W_5__6_), .B(_2923__bF_buf0), .Y(_2210_) );
	OAI21X1 OAI21X1_976 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_4__6_), .C(concatenador_counter_1_bF_buf4), .Y(_2211_) );
	INVX1 INVX1_841 ( .A(micro_hash_synth_1_W_7__6_), .Y(_2212_) );
	AOI21X1 AOI21X1_722 ( .A(concatenador_counter_0_bF_buf13), .B(_2212_), .C(concatenador_counter_1_bF_buf3), .Y(_2213_) );
	OAI21X1 OAI21X1_977 ( .A(concatenador_counter_0_bF_buf12), .B(micro_hash_synth_1_W_6__6_), .C(_2213_), .Y(_2214_) );
	OAI21X1 OAI21X1_978 ( .A(_2210_), .B(_2211_), .C(_2214_), .Y(_2215_) );
	AND2X2 AND2X2_86 ( .A(_2215_), .B(_1633__bF_buf3), .Y(_2216_) );
	AOI21X1 AOI21X1_723 ( .A(concatenador_counter_0_bF_buf11), .B(_3029_), .C(_1657_), .Y(_2217_) );
	OAI21X1 OAI21X1_979 ( .A(concatenador_counter_0_bF_buf10), .B(micro_hash_synth_1_W_0__6_), .C(_2217_), .Y(_2218_) );
	AOI21X1 AOI21X1_724 ( .A(_2923__bF_buf7), .B(_3045_), .C(_1658_), .Y(_2219_) );
	OAI21X1 OAI21X1_980 ( .A(_2923__bF_buf6), .B(micro_hash_synth_1_W_3__6_), .C(_2219_), .Y(_2220_) );
	NAND2X1 NAND2X1_579 ( .A(_2218_), .B(_2220_), .Y(_2221_) );
	OAI21X1 OAI21X1_981 ( .A(_2216_), .B(_2221_), .C(_1643__bF_buf2), .Y(_2222_) );
	NAND2X1 NAND2X1_580 ( .A(_2209_), .B(_2222_), .Y(_2223_) );
	NAND2X1 NAND2X1_581 ( .A(_1680_), .B(_2223_), .Y(_2224_) );
	NAND3X1 NAND3X1_204 ( .A(_2166_), .B(_2194_), .C(_2224_), .Y(_2225_) );
	INVX1 INVX1_842 ( .A(_2225_), .Y(_2226_) );
	AOI21X1 AOI21X1_725 ( .A(_2194_), .B(_2224_), .C(_2166_), .Y(_2227_) );
	OAI21X1 OAI21X1_982 ( .A(_2226_), .B(_2227_), .C(_2162_), .Y(_2228_) );
	INVX1 INVX1_843 ( .A(_2227_), .Y(_2229_) );
	NAND3X1 NAND3X1_205 ( .A(_2161_), .B(_2225_), .C(_2229_), .Y(_2230_) );
	NAND2X1 NAND2X1_582 ( .A(_2228_), .B(_2230_), .Y(_2231_) );
	XNOR2X1 XNOR2X1_37 ( .A(_2160_), .B(_2231_), .Y(_2232_) );
	AOI21X1 AOI21X1_726 ( .A(micro_hash_synth_1_c_6_), .B(_1626_), .C(_1522__bF_buf3), .Y(_2233_) );
	OAI21X1 OAI21X1_983 ( .A(_2232_), .B(_1695_), .C(_2233_), .Y(_1240__6_) );
	NAND2X1 NAND2X1_583 ( .A(_2225_), .B(_2229_), .Y(_2234_) );
	NOR2X1 NOR2X1_419 ( .A(_2161_), .B(_2234_), .Y(_2235_) );
	AOI21X1 AOI21X1_727 ( .A(_2231_), .B(_2160_), .C(_2235_), .Y(_2236_) );
	NOR2X1 NOR2X1_420 ( .A(micro_hash_synth_1_W_21__7_), .B(_2923__bF_buf5), .Y(_2237_) );
	OAI21X1 OAI21X1_984 ( .A(concatenador_counter_0_bF_buf9), .B(micro_hash_synth_1_W_20__7_), .C(concatenador_counter_1_bF_buf2), .Y(_2238_) );
	AOI21X1 AOI21X1_728 ( .A(concatenador_counter_0_bF_buf8), .B(_2959_), .C(concatenador_counter_1_bF_buf1), .Y(_2239_) );
	OAI21X1 OAI21X1_985 ( .A(concatenador_counter_0_bF_buf7), .B(micro_hash_synth_1_W_22__7_), .C(_2239_), .Y(_2240_) );
	OAI21X1 OAI21X1_986 ( .A(_2237_), .B(_2238_), .C(_2240_), .Y(_2241_) );
	INVX1 INVX1_844 ( .A(micro_hash_synth_1_W_18__7_), .Y(_2242_) );
	AOI21X1 AOI21X1_729 ( .A(_2923__bF_buf4), .B(_2242_), .C(_1658_), .Y(_2243_) );
	OAI21X1 OAI21X1_987 ( .A(_2923__bF_buf3), .B(micro_hash_synth_1_W_19__7_), .C(_2243_), .Y(_2244_) );
	NOR2X1 NOR2X1_421 ( .A(micro_hash_synth_1_W_17__7_), .B(_2923__bF_buf2), .Y(_2245_) );
	OAI21X1 OAI21X1_988 ( .A(concatenador_counter_0_bF_buf6), .B(micro_hash_synth_1_W_16__7_), .C(_1630__bF_buf2), .Y(_2246_) );
	OAI21X1 OAI21X1_989 ( .A(_2245_), .B(_2246_), .C(_2244_), .Y(_2247_) );
	AOI21X1 AOI21X1_730 ( .A(_1633__bF_buf2), .B(_2241_), .C(_2247_), .Y(_2248_) );
	NAND2X1 NAND2X1_584 ( .A(_1643__bF_buf1), .B(_2248_), .Y(_2249_) );
	NOR2X1 NOR2X1_422 ( .A(micro_hash_synth_1_W_29__7_), .B(_2923__bF_buf1), .Y(_2250_) );
	OAI21X1 OAI21X1_990 ( .A(concatenador_counter_0_bF_buf5), .B(micro_hash_synth_1_W_28__7_), .C(concatenador_counter_1_bF_buf0), .Y(_2251_) );
	NOR2X1 NOR2X1_423 ( .A(concatenador_counter_0_bF_buf4), .B(micro_hash_synth_1_W_30__7_), .Y(_2252_) );
	OAI21X1 OAI21X1_991 ( .A(_2923__bF_buf0), .B(micro_hash_synth_1_W_31__7_), .C(_1629__bF_buf2), .Y(_2253_) );
	OAI22X1 OAI22X1_296 ( .A(_2250_), .B(_2251_), .C(_2253_), .D(_2252_), .Y(_2254_) );
	NAND2X1 NAND2X1_585 ( .A(_1633__bF_buf1), .B(_2254_), .Y(_2255_) );
	AOI21X1 AOI21X1_731 ( .A(_2923__bF_buf7), .B(_2957_), .C(_1658_), .Y(_2256_) );
	OAI21X1 OAI21X1_992 ( .A(_2923__bF_buf6), .B(micro_hash_synth_1_W_27__7_), .C(_2256_), .Y(_2257_) );
	INVX1 INVX1_845 ( .A(micro_hash_synth_1_W_24__7_), .Y(_2258_) );
	AOI21X1 AOI21X1_732 ( .A(_2923__bF_buf5), .B(_2258_), .C(_1657_), .Y(_2259_) );
	OAI21X1 OAI21X1_993 ( .A(_2923__bF_buf4), .B(micro_hash_synth_1_W_25__7_), .C(_2259_), .Y(_2260_) );
	NAND3X1 NAND3X1_206 ( .A(_2257_), .B(_2260_), .C(_2255_), .Y(_2261_) );
	OAI21X1 OAI21X1_994 ( .A(_1643__bF_buf0), .B(_2261_), .C(_2249_), .Y(_2262_) );
	NAND2X1 NAND2X1_586 ( .A(_1650_), .B(_2262_), .Y(_2263_) );
	NOR2X1 NOR2X1_424 ( .A(micro_hash_synth_1_W_13__7_), .B(_2923__bF_buf3), .Y(_2264_) );
	OAI21X1 OAI21X1_995 ( .A(concatenador_counter_0_bF_buf3), .B(micro_hash_synth_1_W_12__7_), .C(concatenador_counter_1_bF_buf7), .Y(_2265_) );
	INVX1 INVX1_846 ( .A(micro_hash_synth_1_W_15__7_), .Y(_2266_) );
	AOI21X1 AOI21X1_733 ( .A(concatenador_counter_0_bF_buf2), .B(_2266_), .C(concatenador_counter_1_bF_buf6), .Y(_2267_) );
	OAI21X1 OAI21X1_996 ( .A(concatenador_counter_0_bF_buf1), .B(micro_hash_synth_1_W_14__7_), .C(_2267_), .Y(_2268_) );
	OAI21X1 OAI21X1_997 ( .A(_2264_), .B(_2265_), .C(_2268_), .Y(_2269_) );
	AOI21X1 AOI21X1_734 ( .A(_2923__bF_buf2), .B(_3004_), .C(_1657_), .Y(_2270_) );
	OAI21X1 OAI21X1_998 ( .A(_2923__bF_buf1), .B(micro_hash_synth_1_W_9__7_), .C(_2270_), .Y(_2271_) );
	NOR2X1 NOR2X1_425 ( .A(micro_hash_synth_1_W_11__7_), .B(_2923__bF_buf0), .Y(_2272_) );
	OAI21X1 OAI21X1_999 ( .A(concatenador_counter_0_bF_buf0), .B(micro_hash_synth_1_W_10__7_), .C(_1632__bF_buf1), .Y(_2273_) );
	OAI21X1 OAI21X1_1000 ( .A(_2272_), .B(_2273_), .C(_2271_), .Y(_2274_) );
	AOI21X1 AOI21X1_735 ( .A(_1633__bF_buf0), .B(_2269_), .C(_2274_), .Y(_2275_) );
	NAND2X1 NAND2X1_587 ( .A(_1679__bF_buf2), .B(_2275_), .Y(_2276_) );
	NOR2X1 NOR2X1_426 ( .A(micro_hash_synth_1_W_5__7_), .B(_2923__bF_buf7), .Y(_2277_) );
	OAI21X1 OAI21X1_1001 ( .A(concatenador_counter_0_bF_buf13), .B(micro_hash_synth_1_W_4__7_), .C(concatenador_counter_1_bF_buf5), .Y(_2278_) );
	NOR2X1 NOR2X1_427 ( .A(_2278_), .B(_2277_), .Y(_2279_) );
	INVX1 INVX1_847 ( .A(micro_hash_synth_1_W_6__7_), .Y(_2280_) );
	OAI21X1 OAI21X1_1002 ( .A(_2923__bF_buf6), .B(micro_hash_synth_1_W_7__7_), .C(_1629__bF_buf1), .Y(_2281_) );
	AOI21X1 AOI21X1_736 ( .A(_2923__bF_buf5), .B(_2280_), .C(_2281_), .Y(_2282_) );
	OAI21X1 OAI21X1_1003 ( .A(_2282_), .B(_2279_), .C(_1633__bF_buf5), .Y(_2283_) );
	AOI21X1 AOI21X1_737 ( .A(_2923__bF_buf4), .B(_3038_), .C(_1657_), .Y(_2284_) );
	OAI21X1 OAI21X1_1004 ( .A(_2923__bF_buf3), .B(micro_hash_synth_1_W_1__7_), .C(_2284_), .Y(_2285_) );
	AOI21X1 AOI21X1_738 ( .A(_2923__bF_buf2), .B(_3046_), .C(_1658_), .Y(_2286_) );
	OAI21X1 OAI21X1_1005 ( .A(_2923__bF_buf1), .B(micro_hash_synth_1_W_3__7_), .C(_2286_), .Y(_2287_) );
	NAND3X1 NAND3X1_207 ( .A(_2285_), .B(_2287_), .C(_2283_), .Y(_2288_) );
	OAI21X1 OAI21X1_1006 ( .A(_1679__bF_buf1), .B(_2288_), .C(_2276_), .Y(_2289_) );
	NAND2X1 NAND2X1_588 ( .A(_1680_), .B(_2289_), .Y(_2290_) );
	AND2X2 AND2X2_87 ( .A(_2263_), .B(_2290_), .Y(_2291_) );
	XOR2X1 XOR2X1_47 ( .A(micro_hash_synth_1_k_7_), .B(micro_hash_synth_1_x_7_), .Y(_2292_) );
	INVX1 INVX1_848 ( .A(_2292_), .Y(_2293_) );
	NOR2X1 NOR2X1_428 ( .A(_2293_), .B(_2291_), .Y(_2294_) );
	NAND2X1 NAND2X1_589 ( .A(_2263_), .B(_2290_), .Y(_2295_) );
	NOR2X1 NOR2X1_429 ( .A(_2292_), .B(_2295_), .Y(_2296_) );
	OAI22X1 OAI22X1_297 ( .A(_2163_), .B(_2227_), .C(_2294_), .D(_2296_), .Y(_2297_) );
	NOR2X1 NOR2X1_430 ( .A(_2163_), .B(_2227_), .Y(_2298_) );
	NOR2X1 NOR2X1_431 ( .A(_2292_), .B(_2291_), .Y(_2299_) );
	NOR2X1 NOR2X1_432 ( .A(_2293_), .B(_2295_), .Y(_2300_) );
	OAI21X1 OAI21X1_1007 ( .A(_2299_), .B(_2300_), .C(_2298_), .Y(_2301_) );
	NAND2X1 NAND2X1_590 ( .A(_2301_), .B(_2297_), .Y(_2302_) );
	XNOR2X1 XNOR2X1_38 ( .A(_2236_), .B(_2302_), .Y(_2303_) );
	AOI21X1 AOI21X1_739 ( .A(micro_hash_synth_1_c_7_), .B(_1626_), .C(_1522__bF_buf2), .Y(_2304_) );
	OAI21X1 OAI21X1_1008 ( .A(_2303_), .B(_1695_), .C(_2304_), .Y(_1240__7_) );
	OAI21X1 OAI21X1_1009 ( .A(_1512_), .B(_1614__bF_buf2), .C(_1523__bF_buf3), .Y(_1239__0_) );
	NOR2X1 NOR2X1_433 ( .A(_1515_), .B(_1616_), .Y(_1239__1_) );
	INVX1 INVX1_849 ( .A(micro_hash_synth_1_b_2_), .Y(_2305_) );
	NOR2X1 NOR2X1_434 ( .A(_2305_), .B(_1616_), .Y(_1239__2_) );
	OAI21X1 OAI21X1_1010 ( .A(_1533_), .B(_1614__bF_buf1), .C(_1523__bF_buf2), .Y(_1239__3_) );
	OAI21X1 OAI21X1_1011 ( .A(micro_hash_synth_1_b_4_), .B(_1614__bF_buf0), .C(_1523__bF_buf1), .Y(_2306_) );
	AOI21X1 AOI21X1_740 ( .A(_1628_), .B(_1793_), .C(_2306_), .Y(_1239__4_) );
	INVX1 INVX1_850 ( .A(micro_hash_synth_1_c_1_), .Y(_2307_) );
	OAI21X1 OAI21X1_1012 ( .A(micro_hash_synth_1_b_5_), .B(_1614__bF_buf3), .C(_1523__bF_buf0), .Y(_2308_) );
	AOI21X1 AOI21X1_741 ( .A(_2307_), .B(_1793_), .C(_2308_), .Y(_1239__5_) );
	INVX1 INVX1_851 ( .A(micro_hash_synth_1_c_2_), .Y(_2309_) );
	OAI21X1 OAI21X1_1013 ( .A(micro_hash_synth_1_b_6_), .B(_1614__bF_buf2), .C(_1523__bF_buf3), .Y(_2310_) );
	AOI21X1 AOI21X1_742 ( .A(_2309_), .B(_1793_), .C(_2310_), .Y(_1239__6_) );
	INVX1 INVX1_852 ( .A(micro_hash_synth_1_b_7_), .Y(_2311_) );
	NOR2X1 NOR2X1_435 ( .A(micro_hash_synth_1_c_3_), .B(_1626_), .Y(_2312_) );
	AOI22X1 AOI22X1_35 ( .A(_2311_), .B(_1615_), .C(_2312_), .D(_1523__bF_buf2), .Y(_1239__7_) );
	XNOR2X1 XNOR2X1_39 ( .A(micro_hash_synth_1_b_0_), .B(micro_hash_synth_1_c_0_), .Y(_2313_) );
	AOI21X1 AOI21X1_743 ( .A(micro_hash_synth_1_a_0_), .B(_1626_), .C(_1522__bF_buf1), .Y(_2314_) );
	OAI21X1 OAI21X1_1014 ( .A(_1695_), .B(_2313_), .C(_2314_), .Y(_1238__0_) );
	NOR2X1 NOR2X1_436 ( .A(micro_hash_synth_1_b_1_), .B(_2307_), .Y(_2315_) );
	NOR2X1 NOR2X1_437 ( .A(micro_hash_synth_1_c_1_), .B(_1515_), .Y(_2316_) );
	OAI21X1 OAI21X1_1015 ( .A(_2315_), .B(_2316_), .C(_1793_), .Y(_2317_) );
	OAI22X1 OAI22X1_298 ( .A(_1568_), .B(_1616_), .C(_2317_), .D(_3022__bF_buf5), .Y(_1238__1_) );
	INVX1 INVX1_853 ( .A(micro_hash_synth_1_a_2_), .Y(_2318_) );
	NOR2X1 NOR2X1_438 ( .A(micro_hash_synth_1_b_2_), .B(_2309_), .Y(_2319_) );
	NOR2X1 NOR2X1_439 ( .A(micro_hash_synth_1_c_2_), .B(_2305_), .Y(_2320_) );
	OAI21X1 OAI21X1_1016 ( .A(_2319_), .B(_2320_), .C(_1793_), .Y(_2321_) );
	OAI22X1 OAI22X1_299 ( .A(_2318_), .B(_1616_), .C(_2321_), .D(_3022__bF_buf4), .Y(_1238__2_) );
	NAND2X1 NAND2X1_591 ( .A(micro_hash_synth_1_a_3_), .B(_1615_), .Y(_2322_) );
	INVX1 INVX1_854 ( .A(micro_hash_synth_1_c_3_), .Y(_2323_) );
	NOR2X1 NOR2X1_440 ( .A(micro_hash_synth_1_b_3_), .B(_2323_), .Y(_2324_) );
	NOR2X1 NOR2X1_441 ( .A(micro_hash_synth_1_c_3_), .B(_1533_), .Y(_2325_) );
	OAI21X1 OAI21X1_1017 ( .A(_2324_), .B(_2325_), .C(_1793_), .Y(_2326_) );
	OAI21X1 OAI21X1_1018 ( .A(_2326_), .B(_3022__bF_buf3), .C(_2322_), .Y(_1238__3_) );
	INVX1 INVX1_855 ( .A(micro_hash_synth_1_a_4_), .Y(_2327_) );
	INVX1 INVX1_856 ( .A(micro_hash_synth_1_c_4_), .Y(_2328_) );
	NOR2X1 NOR2X1_442 ( .A(micro_hash_synth_1_b_4_), .B(_2328_), .Y(_2329_) );
	INVX1 INVX1_857 ( .A(micro_hash_synth_1_b_4_), .Y(_2330_) );
	NOR2X1 NOR2X1_443 ( .A(micro_hash_synth_1_c_4_), .B(_2330_), .Y(_2331_) );
	OAI21X1 OAI21X1_1019 ( .A(_2329_), .B(_2331_), .C(_1793_), .Y(_2332_) );
	OAI22X1 OAI22X1_300 ( .A(_2327_), .B(_1616_), .C(_2332_), .D(_3022__bF_buf2), .Y(_1238__4_) );
	NAND2X1 NAND2X1_592 ( .A(micro_hash_synth_1_a_5_), .B(_1615_), .Y(_2333_) );
	INVX1 INVX1_858 ( .A(micro_hash_synth_1_c_5_), .Y(_2334_) );
	NOR2X1 NOR2X1_444 ( .A(micro_hash_synth_1_b_5_), .B(_2334_), .Y(_2335_) );
	AND2X2 AND2X2_88 ( .A(_2334_), .B(micro_hash_synth_1_b_5_), .Y(_2336_) );
	OAI21X1 OAI21X1_1020 ( .A(_2335_), .B(_2336_), .C(_1793_), .Y(_2337_) );
	OAI21X1 OAI21X1_1021 ( .A(_2337_), .B(_3022__bF_buf1), .C(_2333_), .Y(_1238__5_) );
	INVX1 INVX1_859 ( .A(micro_hash_synth_1_c_6_), .Y(_2338_) );
	NOR2X1 NOR2X1_445 ( .A(micro_hash_synth_1_b_6_), .B(_2338_), .Y(_2339_) );
	AND2X2 AND2X2_89 ( .A(_2338_), .B(micro_hash_synth_1_b_6_), .Y(_2340_) );
	OAI21X1 OAI21X1_1022 ( .A(_2339_), .B(_2340_), .C(_1793_), .Y(_2341_) );
	OAI22X1 OAI22X1_301 ( .A(_1608_), .B(_1616_), .C(_2341_), .D(_3022__bF_buf0), .Y(_1238__6_) );
	INVX1 INVX1_860 ( .A(micro_hash_synth_1_a_7_), .Y(_2342_) );
	AND2X2 AND2X2_90 ( .A(_2311_), .B(micro_hash_synth_1_c_7_), .Y(_2343_) );
	NOR2X1 NOR2X1_446 ( .A(micro_hash_synth_1_c_7_), .B(_2311_), .Y(_2344_) );
	OAI21X1 OAI21X1_1023 ( .A(_2343_), .B(_2344_), .C(_1793_), .Y(_2345_) );
	OAI22X1 OAI22X1_302 ( .A(_2342_), .B(_1616_), .C(_2345_), .D(_3022__bF_buf5), .Y(_1238__7_) );
	XNOR2X1 XNOR2X1_40 ( .A(micro_hash_synth_1_c_0_), .B(Hhash_synth1_16_), .Y(_2346_) );
	NAND2X1 NAND2X1_593 ( .A(Hhash_synth1_16_), .B(_1523__bF_buf1), .Y(_2347_) );
	AOI22X1 AOI22X1_36 ( .A(_1506__bF_buf3), .B(_2346_), .C(_1510_), .D(_2347_), .Y(_1237__16_) );
	INVX1 INVX1_861 ( .A(Hhash_synth1_17_), .Y(_2348_) );
	NOR2X1 NOR2X1_447 ( .A(_2307_), .B(_2348_), .Y(_2349_) );
	NOR2X1 NOR2X1_448 ( .A(micro_hash_synth_1_c_1_), .B(Hhash_synth1_17_), .Y(_2350_) );
	NOR2X1 NOR2X1_449 ( .A(_2350_), .B(_2349_), .Y(_2351_) );
	NAND3X1 NAND3X1_208 ( .A(micro_hash_synth_1_c_0_), .B(Hhash_synth1_16_), .C(_2351_), .Y(_2352_) );
	NAND2X1 NAND2X1_594 ( .A(micro_hash_synth_1_c_0_), .B(Hhash_synth1_16_), .Y(_2353_) );
	OAI21X1 OAI21X1_1024 ( .A(_2349_), .B(_2350_), .C(_2353_), .Y(_2354_) );
	NAND3X1 NAND3X1_209 ( .A(_2352_), .B(_2354_), .C(_1506__bF_buf2), .Y(_2355_) );
	OAI21X1 OAI21X1_1025 ( .A(_2928_), .B(Hhash_synth1_17_), .C(_1507_), .Y(_2356_) );
	NAND3X1 NAND3X1_210 ( .A(reset_L_bF_buf1), .B(_2355_), .C(_2356_), .Y(_1237__17_) );
	OAI21X1 OAI21X1_1026 ( .A(Hhash_synth1_18_), .B(_1522__bF_buf0), .C(_1510_), .Y(_2357_) );
	OAI21X1 OAI21X1_1027 ( .A(_2307_), .B(_2348_), .C(_2352_), .Y(_2358_) );
	INVX1 INVX1_862 ( .A(Hhash_synth1_18_), .Y(_2359_) );
	NOR2X1 NOR2X1_450 ( .A(_2309_), .B(_2359_), .Y(_2360_) );
	NOR2X1 NOR2X1_451 ( .A(micro_hash_synth_1_c_2_), .B(Hhash_synth1_18_), .Y(_2361_) );
	NOR2X1 NOR2X1_452 ( .A(_2361_), .B(_2360_), .Y(_2362_) );
	NOR2X1 NOR2X1_453 ( .A(_2362_), .B(_2358_), .Y(_2363_) );
	NAND2X1 NAND2X1_595 ( .A(_2362_), .B(_2358_), .Y(_2364_) );
	NAND2X1 NAND2X1_596 ( .A(_2364_), .B(_1506__bF_buf1), .Y(_2365_) );
	OAI21X1 OAI21X1_1028 ( .A(_2365_), .B(_2363_), .C(_2357_), .Y(_1237__18_) );
	AOI21X1 AOI21X1_744 ( .A(_2362_), .B(_2358_), .C(_2360_), .Y(_2366_) );
	INVX1 INVX1_863 ( .A(Hhash_synth1_19_), .Y(_2367_) );
	NOR2X1 NOR2X1_454 ( .A(_2323_), .B(_2367_), .Y(_2368_) );
	NOR2X1 NOR2X1_455 ( .A(micro_hash_synth_1_c_3_), .B(Hhash_synth1_19_), .Y(_2369_) );
	NOR2X1 NOR2X1_456 ( .A(_2369_), .B(_2368_), .Y(_2370_) );
	XOR2X1 XOR2X1_48 ( .A(_2366_), .B(_2370_), .Y(_2371_) );
	OAI21X1 OAI21X1_1029 ( .A(Hhash_synth1_19_), .B(_1522__bF_buf3), .C(_1510_), .Y(_2372_) );
	OAI21X1 OAI21X1_1030 ( .A(_1507_), .B(_2371_), .C(_2372_), .Y(_1237__19_) );
	XOR2X1 XOR2X1_49 ( .A(micro_hash_synth_1_c_4_), .B(Hhash_synth1_20_), .Y(_2373_) );
	INVX1 INVX1_864 ( .A(_2373_), .Y(_2374_) );
	OAI21X1 OAI21X1_1031 ( .A(_2323_), .B(_2367_), .C(_2366_), .Y(_2375_) );
	OAI21X1 OAI21X1_1032 ( .A(micro_hash_synth_1_c_3_), .B(Hhash_synth1_19_), .C(_2375_), .Y(_2376_) );
	NAND2X1 NAND2X1_597 ( .A(_2374_), .B(_2376_), .Y(_2377_) );
	NOR2X1 NOR2X1_457 ( .A(_2374_), .B(_2376_), .Y(_2378_) );
	INVX1 INVX1_865 ( .A(_2378_), .Y(_2379_) );
	NAND2X1 NAND2X1_598 ( .A(_2377_), .B(_2379_), .Y(_2380_) );
	OAI21X1 OAI21X1_1033 ( .A(Hhash_synth1_20_), .B(_1522__bF_buf2), .C(_1510_), .Y(_2381_) );
	OAI21X1 OAI21X1_1034 ( .A(_2380_), .B(_1507_), .C(_2381_), .Y(_1237__20_) );
	OAI21X1 OAI21X1_1035 ( .A(Hhash_synth1_21_), .B(_1522__bF_buf1), .C(_1510_), .Y(_2382_) );
	AOI21X1 AOI21X1_745 ( .A(micro_hash_synth_1_c_4_), .B(Hhash_synth1_20_), .C(_2378_), .Y(_2383_) );
	INVX1 INVX1_866 ( .A(Hhash_synth1_21_), .Y(_2384_) );
	NOR2X1 NOR2X1_458 ( .A(_2334_), .B(_2384_), .Y(_2385_) );
	NOR2X1 NOR2X1_459 ( .A(micro_hash_synth_1_c_5_), .B(Hhash_synth1_21_), .Y(_2386_) );
	NOR2X1 NOR2X1_460 ( .A(_2386_), .B(_2385_), .Y(_2387_) );
	XOR2X1 XOR2X1_50 ( .A(_2383_), .B(_2387_), .Y(_2388_) );
	OAI21X1 OAI21X1_1036 ( .A(_2388_), .B(_1507_), .C(_2382_), .Y(_1237__21_) );
	OAI21X1 OAI21X1_1037 ( .A(Hhash_synth1_22_), .B(_1522__bF_buf0), .C(_1510_), .Y(_2389_) );
	XOR2X1 XOR2X1_51 ( .A(micro_hash_synth_1_c_6_), .B(Hhash_synth1_22_), .Y(_2390_) );
	INVX1 INVX1_867 ( .A(_2385_), .Y(_2391_) );
	OAI21X1 OAI21X1_1038 ( .A(_2383_), .B(_2386_), .C(_2391_), .Y(_2392_) );
	NOR2X1 NOR2X1_461 ( .A(_2390_), .B(_2392_), .Y(_2393_) );
	NAND2X1 NAND2X1_599 ( .A(_2390_), .B(_2392_), .Y(_2394_) );
	NAND2X1 NAND2X1_600 ( .A(_1506__bF_buf0), .B(_2394_), .Y(_2395_) );
	OAI21X1 OAI21X1_1039 ( .A(_2395_), .B(_2393_), .C(_2389_), .Y(_1237__22_) );
	OAI21X1 OAI21X1_1040 ( .A(Hhash_synth1_23_), .B(_1522__bF_buf3), .C(_1510_), .Y(_2396_) );
	INVX1 INVX1_868 ( .A(Hhash_synth1_22_), .Y(_2397_) );
	OAI21X1 OAI21X1_1041 ( .A(_2338_), .B(_2397_), .C(_2394_), .Y(_2398_) );
	XNOR2X1 XNOR2X1_41 ( .A(micro_hash_synth_1_c_7_), .B(Hhash_synth1_23_), .Y(_2399_) );
	INVX1 INVX1_869 ( .A(_2399_), .Y(_2400_) );
	AND2X2 AND2X2_91 ( .A(_2398_), .B(_2400_), .Y(_2401_) );
	OAI21X1 OAI21X1_1042 ( .A(_2398_), .B(_2400_), .C(_1506__bF_buf3), .Y(_2402_) );
	OAI21X1 OAI21X1_1043 ( .A(_2401_), .B(_2402_), .C(_2396_), .Y(_1237__23_) );
	NAND3X1 NAND3X1_211 ( .A(_1512_), .B(_1565_), .C(_1614__bF_buf1), .Y(_2403_) );
	OAI21X1 OAI21X1_1044 ( .A(micro_hash_synth_1_x_0_), .B(_1614__bF_buf0), .C(_2403_), .Y(_2404_) );
	XNOR2X1 XNOR2X1_42 ( .A(micro_hash_synth_1_b_0_), .B(micro_hash_synth_1_a_0_), .Y(_2405_) );
	NAND2X1 NAND2X1_601 ( .A(_1622_), .B(_1523__bF_buf0), .Y(_2406_) );
	OAI22X1 OAI22X1_303 ( .A(_2405_), .B(_2406_), .C(_2404_), .D(_1627_), .Y(_1243__0_) );
	NAND3X1 NAND3X1_212 ( .A(_1515_), .B(_1568_), .C(_1614__bF_buf3), .Y(_2407_) );
	OAI21X1 OAI21X1_1045 ( .A(micro_hash_synth_1_x_1_), .B(_1614__bF_buf2), .C(_2407_), .Y(_2408_) );
	XNOR2X1 XNOR2X1_43 ( .A(micro_hash_synth_1_b_1_), .B(micro_hash_synth_1_a_1_), .Y(_2409_) );
	OAI22X1 OAI22X1_304 ( .A(_2406_), .B(_2409_), .C(_2408_), .D(_1627_), .Y(_1243__1_) );
	NAND3X1 NAND3X1_213 ( .A(_2305_), .B(_2318_), .C(_1614__bF_buf1), .Y(_2410_) );
	OAI21X1 OAI21X1_1046 ( .A(micro_hash_synth_1_x_2_), .B(_1614__bF_buf0), .C(_2410_), .Y(_2411_) );
	XNOR2X1 XNOR2X1_44 ( .A(micro_hash_synth_1_b_2_), .B(micro_hash_synth_1_a_2_), .Y(_2412_) );
	OAI22X1 OAI22X1_305 ( .A(_2406_), .B(_2412_), .C(_2411_), .D(_1627_), .Y(_1243__2_) );
	XOR2X1 XOR2X1_52 ( .A(micro_hash_synth_1_b_3_), .B(micro_hash_synth_1_a_3_), .Y(_2413_) );
	OAI21X1 OAI21X1_1047 ( .A(_1522__bF_buf2), .B(_2413_), .C(_1627_), .Y(_2414_) );
	OAI21X1 OAI21X1_1048 ( .A(micro_hash_synth_1_b_3_), .B(micro_hash_synth_1_a_3_), .C(_1614__bF_buf3), .Y(_2415_) );
	OAI21X1 OAI21X1_1049 ( .A(_1909_), .B(_1614__bF_buf2), .C(_2415_), .Y(_2416_) );
	NAND2X1 NAND2X1_602 ( .A(_1621_), .B(_2416_), .Y(_2417_) );
	NAND2X1 NAND2X1_603 ( .A(_2414_), .B(_2417_), .Y(_1243__3_) );
	NAND3X1 NAND3X1_214 ( .A(_2330_), .B(_2327_), .C(_1614__bF_buf1), .Y(_2418_) );
	OAI21X1 OAI21X1_1050 ( .A(micro_hash_synth_1_x_4_), .B(_1614__bF_buf0), .C(_2418_), .Y(_2419_) );
	XNOR2X1 XNOR2X1_45 ( .A(micro_hash_synth_1_b_4_), .B(micro_hash_synth_1_a_4_), .Y(_2420_) );
	OAI22X1 OAI22X1_306 ( .A(_2406_), .B(_2420_), .C(_2419_), .D(_1627_), .Y(_1243__4_) );
	NOR2X1 NOR2X1_462 ( .A(micro_hash_synth_1_b_5_), .B(micro_hash_synth_1_a_5_), .Y(_2421_) );
	OAI21X1 OAI21X1_1051 ( .A(_1501_), .B(_1503_), .C(_2421_), .Y(_2422_) );
	OAI21X1 OAI21X1_1052 ( .A(micro_hash_synth_1_x_5_), .B(_1614__bF_buf3), .C(_2422_), .Y(_2423_) );
	XNOR2X1 XNOR2X1_46 ( .A(micro_hash_synth_1_b_5_), .B(micro_hash_synth_1_a_5_), .Y(_2424_) );
	OAI22X1 OAI22X1_307 ( .A(_2406_), .B(_2424_), .C(_2423_), .D(_1627_), .Y(_1243__5_) );
	NOR2X1 NOR2X1_463 ( .A(micro_hash_synth_1_b_6_), .B(micro_hash_synth_1_a_6_), .Y(_2425_) );
	OAI21X1 OAI21X1_1053 ( .A(_1501_), .B(_1503_), .C(_2425_), .Y(_2426_) );
	OAI21X1 OAI21X1_1054 ( .A(micro_hash_synth_1_x_6_), .B(_1614__bF_buf2), .C(_2426_), .Y(_2427_) );
	XNOR2X1 XNOR2X1_47 ( .A(micro_hash_synth_1_b_6_), .B(micro_hash_synth_1_a_6_), .Y(_2428_) );
	OAI22X1 OAI22X1_308 ( .A(_2406_), .B(_2428_), .C(_2427_), .D(_1627_), .Y(_1243__6_) );
	XOR2X1 XOR2X1_53 ( .A(micro_hash_synth_1_b_7_), .B(micro_hash_synth_1_a_7_), .Y(_2429_) );
	OAI21X1 OAI21X1_1055 ( .A(_1522__bF_buf1), .B(_2429_), .C(_1627_), .Y(_2430_) );
	NAND2X1 NAND2X1_604 ( .A(_2311_), .B(_2342_), .Y(_2431_) );
	NOR2X1 NOR2X1_464 ( .A(_2431_), .B(_1626_), .Y(_2432_) );
	OAI21X1 OAI21X1_1056 ( .A(_1614__bF_buf1), .B(micro_hash_synth_1_x_7_), .C(_1621_), .Y(_2433_) );
	OAI21X1 OAI21X1_1057 ( .A(_2433_), .B(_2432_), .C(_2430_), .Y(_1243__7_) );
	INVX1 INVX1_870 ( .A(micro_hash_synth_1_W_24__0_), .Y(_2434_) );
	XOR2X1 XOR2X1_54 ( .A(micro_hash_synth_1_W_10__0_), .B(micro_hash_synth_1_W_15__0_), .Y(_2435_) );
	NOR2X1 NOR2X1_465 ( .A(micro_hash_synth_1_W_21__0_), .B(_2435_), .Y(_2436_) );
	OAI22X1 OAI22X1_309 ( .A(_2925__bF_buf15), .B(_2436_), .C(_2930__bF_buf9), .D(_2434_), .Y(_1406_) );
	INVX1 INVX1_871 ( .A(micro_hash_synth_1_W_21__1_), .Y(_2437_) );
	OAI21X1 OAI21X1_1058 ( .A(_1736_), .B(micro_hash_synth_1_W_15__1_), .C(_2437_), .Y(_2438_) );
	AOI21X1 AOI21X1_746 ( .A(_1736_), .B(micro_hash_synth_1_W_15__1_), .C(_2438_), .Y(_2439_) );
	OAI22X1 OAI22X1_310 ( .A(_2925__bF_buf14), .B(_2439_), .C(_2930__bF_buf8), .D(_1723_), .Y(_1407_) );
	INVX1 INVX1_872 ( .A(micro_hash_synth_1_W_21__2_), .Y(_2440_) );
	OAI21X1 OAI21X1_1059 ( .A(_1836_), .B(micro_hash_synth_1_W_15__2_), .C(_2440_), .Y(_2441_) );
	AOI21X1 AOI21X1_747 ( .A(_1836_), .B(micro_hash_synth_1_W_15__2_), .C(_2441_), .Y(_2442_) );
	OAI22X1 OAI22X1_311 ( .A(_2925__bF_buf13), .B(_2442_), .C(_2930__bF_buf7), .D(_1819_), .Y(_1408_) );
	INVX1 INVX1_873 ( .A(micro_hash_synth_1_W_21__3_), .Y(_2443_) );
	OAI21X1 OAI21X1_1060 ( .A(_1951_), .B(micro_hash_synth_1_W_15__3_), .C(_2443_), .Y(_2444_) );
	AOI21X1 AOI21X1_748 ( .A(_1951_), .B(micro_hash_synth_1_W_15__3_), .C(_2444_), .Y(_2445_) );
	OAI22X1 OAI22X1_312 ( .A(_2925__bF_buf12), .B(_2445_), .C(_2930__bF_buf6), .D(_1919_), .Y(_1409_) );
	INVX1 INVX1_874 ( .A(micro_hash_synth_1_W_21__4_), .Y(_2446_) );
	OAI21X1 OAI21X1_1061 ( .A(_2017_), .B(micro_hash_synth_1_W_15__4_), .C(_2446_), .Y(_2447_) );
	AOI21X1 AOI21X1_749 ( .A(_2017_), .B(micro_hash_synth_1_W_15__4_), .C(_2447_), .Y(_2448_) );
	OAI22X1 OAI22X1_313 ( .A(_2925__bF_buf11), .B(_2448_), .C(_2930__bF_buf5), .D(_2003_), .Y(_1410_) );
	INVX1 INVX1_875 ( .A(micro_hash_synth_1_W_21__5_), .Y(_2449_) );
	OAI21X1 OAI21X1_1062 ( .A(_2119_), .B(micro_hash_synth_1_W_15__5_), .C(_2449_), .Y(_2450_) );
	AOI21X1 AOI21X1_750 ( .A(_2119_), .B(micro_hash_synth_1_W_15__5_), .C(_2450_), .Y(_2451_) );
	OAI22X1 OAI22X1_314 ( .A(_2925__bF_buf10), .B(_2451_), .C(_2930__bF_buf4), .D(_2105_), .Y(_1411_) );
	INVX1 INVX1_876 ( .A(micro_hash_synth_1_W_21__6_), .Y(_2452_) );
	OAI21X1 OAI21X1_1063 ( .A(_2205_), .B(micro_hash_synth_1_W_15__6_), .C(_2452_), .Y(_2453_) );
	AOI21X1 AOI21X1_751 ( .A(_2205_), .B(micro_hash_synth_1_W_15__6_), .C(_2453_), .Y(_2454_) );
	OAI22X1 OAI22X1_315 ( .A(_2925__bF_buf9), .B(_2454_), .C(_2930__bF_buf3), .D(_2186_), .Y(_1413_) );
	INVX1 INVX1_877 ( .A(micro_hash_synth_1_W_10__7_), .Y(_2455_) );
	INVX1 INVX1_878 ( .A(micro_hash_synth_1_W_21__7_), .Y(_2456_) );
	OAI21X1 OAI21X1_1064 ( .A(_2455_), .B(micro_hash_synth_1_W_15__7_), .C(_2456_), .Y(_2457_) );
	AOI21X1 AOI21X1_752 ( .A(_2455_), .B(micro_hash_synth_1_W_15__7_), .C(_2457_), .Y(_2458_) );
	OAI22X1 OAI22X1_316 ( .A(_2925__bF_buf8), .B(_2458_), .C(_2930__bF_buf2), .D(_2258_), .Y(_1414_) );
	INVX8 INVX8_8 ( .A(_2930__bF_buf1), .Y(_2459_) );
	NAND2X1 NAND2X1_605 ( .A(micro_hash_synth_1_W_23__0_), .B(_2459__bF_buf6), .Y(_2460_) );
	XOR2X1 XOR2X1_55 ( .A(micro_hash_synth_1_W_9__0_), .B(micro_hash_synth_1_W_14__0_), .Y(_2461_) );
	NOR2X1 NOR2X1_466 ( .A(micro_hash_synth_1_W_20__0_), .B(_2461_), .Y(_2462_) );
	OAI21X1 OAI21X1_1065 ( .A(_2925__bF_buf7), .B(_2462_), .C(_2460_), .Y(_1415_) );
	XOR2X1 XOR2X1_56 ( .A(micro_hash_synth_1_W_9__1_), .B(micro_hash_synth_1_W_14__1_), .Y(_2463_) );
	NOR2X1 NOR2X1_467 ( .A(micro_hash_synth_1_W_20__1_), .B(_2463_), .Y(_2464_) );
	OAI22X1 OAI22X1_317 ( .A(_2925__bF_buf6), .B(_2464_), .C(_2930__bF_buf0), .D(_2935_), .Y(_1416_) );
	XOR2X1 XOR2X1_57 ( .A(micro_hash_synth_1_W_9__2_), .B(micro_hash_synth_1_W_14__2_), .Y(_2465_) );
	NOR2X1 NOR2X1_468 ( .A(micro_hash_synth_1_W_20__2_), .B(_2465_), .Y(_2466_) );
	OAI22X1 OAI22X1_318 ( .A(_2925__bF_buf5), .B(_2466_), .C(_2930__bF_buf13), .D(_2940_), .Y(_1417_) );
	NAND2X1 NAND2X1_606 ( .A(micro_hash_synth_1_W_23__3_), .B(_2459__bF_buf5), .Y(_2467_) );
	XOR2X1 XOR2X1_58 ( .A(micro_hash_synth_1_W_9__3_), .B(micro_hash_synth_1_W_14__3_), .Y(_2468_) );
	NOR2X1 NOR2X1_469 ( .A(micro_hash_synth_1_W_20__3_), .B(_2468_), .Y(_2469_) );
	OAI21X1 OAI21X1_1066 ( .A(_2925__bF_buf4), .B(_2469_), .C(_2467_), .Y(_1418_) );
	NAND2X1 NAND2X1_607 ( .A(micro_hash_synth_1_W_23__4_), .B(_2459__bF_buf4), .Y(_2470_) );
	XOR2X1 XOR2X1_59 ( .A(micro_hash_synth_1_W_9__4_), .B(micro_hash_synth_1_W_14__4_), .Y(_2471_) );
	NOR2X1 NOR2X1_470 ( .A(micro_hash_synth_1_W_20__4_), .B(_2471_), .Y(_2472_) );
	OAI21X1 OAI21X1_1067 ( .A(_2925__bF_buf3), .B(_2472_), .C(_2470_), .Y(_1419_) );
	NAND2X1 NAND2X1_608 ( .A(micro_hash_synth_1_W_23__5_), .B(_2459__bF_buf3), .Y(_2473_) );
	XOR2X1 XOR2X1_60 ( .A(micro_hash_synth_1_W_9__5_), .B(micro_hash_synth_1_W_14__5_), .Y(_2474_) );
	NOR2X1 NOR2X1_471 ( .A(micro_hash_synth_1_W_20__5_), .B(_2474_), .Y(_2475_) );
	OAI21X1 OAI21X1_1068 ( .A(_2925__bF_buf2), .B(_2475_), .C(_2473_), .Y(_1420_) );
	INVX1 INVX1_879 ( .A(micro_hash_synth_1_W_20__6_), .Y(_2476_) );
	OAI21X1 OAI21X1_1069 ( .A(_2202_), .B(micro_hash_synth_1_W_14__6_), .C(_2476_), .Y(_2477_) );
	AOI21X1 AOI21X1_753 ( .A(_2202_), .B(micro_hash_synth_1_W_14__6_), .C(_2477_), .Y(_2478_) );
	OAI22X1 OAI22X1_319 ( .A(_2925__bF_buf1), .B(_2478_), .C(_2930__bF_buf12), .D(_2954_), .Y(_1421_) );
	XOR2X1 XOR2X1_61 ( .A(micro_hash_synth_1_W_9__7_), .B(micro_hash_synth_1_W_14__7_), .Y(_2479_) );
	NOR2X1 NOR2X1_472 ( .A(micro_hash_synth_1_W_20__7_), .B(_2479_), .Y(_2480_) );
	OAI22X1 OAI22X1_320 ( .A(_2925__bF_buf0), .B(_2480_), .C(_2930__bF_buf11), .D(_2959_), .Y(_1422_) );
	INVX1 INVX1_880 ( .A(micro_hash_synth_1_W_7__0_), .Y(_2481_) );
	INVX1 INVX1_881 ( .A(bloque_in_56_), .Y(_2482_) );
	OAI22X1 OAI22X1_321 ( .A(_2482_), .B(_2925__bF_buf15), .C(_2930__bF_buf10), .D(_2481_), .Y(_1424_) );
	INVX1 INVX1_882 ( .A(bloque_in_57_), .Y(_2483_) );
	OAI22X1 OAI22X1_322 ( .A(_2483_), .B(_2925__bF_buf14), .C(_2930__bF_buf9), .D(_1750_), .Y(_1425_) );
	INVX1 INVX1_883 ( .A(bloque_in_58_), .Y(_2484_) );
	OAI22X1 OAI22X1_323 ( .A(_2484_), .B(_2925__bF_buf13), .C(_2930__bF_buf8), .D(_1884_), .Y(_1426_) );
	INVX1 INVX1_884 ( .A(micro_hash_synth_1_W_7__3_), .Y(_2485_) );
	INVX1 INVX1_885 ( .A(bloque_in_59_), .Y(_2486_) );
	OAI22X1 OAI22X1_324 ( .A(_2486_), .B(_2925__bF_buf12), .C(_2930__bF_buf7), .D(_2485_), .Y(_1427_) );
	INVX1 INVX1_886 ( .A(micro_hash_synth_1_W_7__4_), .Y(_2487_) );
	INVX1 INVX1_887 ( .A(bloque_in_60_), .Y(_2488_) );
	OAI22X1 OAI22X1_325 ( .A(_2488_), .B(_2925__bF_buf11), .C(_2930__bF_buf6), .D(_2487_), .Y(_1428_) );
	INVX1 INVX1_888 ( .A(micro_hash_synth_1_W_7__5_), .Y(_2489_) );
	INVX1 INVX1_889 ( .A(bloque_in_61_), .Y(_2490_) );
	OAI22X1 OAI22X1_326 ( .A(_2490_), .B(_2925__bF_buf10), .C(_2930__bF_buf5), .D(_2489_), .Y(_1429_) );
	INVX1 INVX1_890 ( .A(bloque_in_62_), .Y(_2491_) );
	OAI22X1 OAI22X1_327 ( .A(_2491_), .B(_2925__bF_buf9), .C(_2930__bF_buf4), .D(_2212_), .Y(_1430_) );
	INVX1 INVX1_891 ( .A(micro_hash_synth_1_W_7__7_), .Y(_2492_) );
	INVX1 INVX1_892 ( .A(bloque_in_63_), .Y(_2493_) );
	OAI22X1 OAI22X1_328 ( .A(_2493_), .B(_2925__bF_buf8), .C(_2930__bF_buf3), .D(_2492_), .Y(_1431_) );
	NAND2X1 NAND2X1_609 ( .A(micro_hash_synth_1_W_22__0_), .B(_2459__bF_buf2), .Y(_2494_) );
	INVX1 INVX1_893 ( .A(micro_hash_synth_1_W_19__0_), .Y(_2495_) );
	OAI21X1 OAI21X1_1070 ( .A(_2990_), .B(micro_hash_synth_1_W_13__0_), .C(_2495_), .Y(_2496_) );
	AOI21X1 AOI21X1_754 ( .A(_2990_), .B(micro_hash_synth_1_W_13__0_), .C(_2496_), .Y(_2497_) );
	OAI21X1 OAI21X1_1071 ( .A(_2925__bF_buf7), .B(_2497_), .C(_2494_), .Y(_1432_) );
	INVX1 INVX1_894 ( .A(micro_hash_synth_1_W_19__1_), .Y(_2498_) );
	OAI21X1 OAI21X1_1072 ( .A(_2992_), .B(micro_hash_synth_1_W_13__1_), .C(_2498_), .Y(_2499_) );
	AOI21X1 AOI21X1_755 ( .A(_2992_), .B(micro_hash_synth_1_W_13__1_), .C(_2499_), .Y(_2500_) );
	OAI22X1 OAI22X1_329 ( .A(_2925__bF_buf6), .B(_2500_), .C(_2930__bF_buf2), .D(_2967_), .Y(_1433_) );
	INVX1 INVX1_895 ( .A(micro_hash_synth_1_W_19__2_), .Y(_2501_) );
	OAI21X1 OAI21X1_1073 ( .A(_2994_), .B(micro_hash_synth_1_W_13__2_), .C(_2501_), .Y(_2502_) );
	AOI21X1 AOI21X1_756 ( .A(_2994_), .B(micro_hash_synth_1_W_13__2_), .C(_2502_), .Y(_2503_) );
	OAI22X1 OAI22X1_330 ( .A(_2925__bF_buf5), .B(_2503_), .C(_2930__bF_buf1), .D(_2972_), .Y(_1435_) );
	NAND2X1 NAND2X1_610 ( .A(micro_hash_synth_1_W_22__3_), .B(_2459__bF_buf1), .Y(_2504_) );
	INVX1 INVX1_896 ( .A(micro_hash_synth_1_W_19__3_), .Y(_2505_) );
	OAI21X1 OAI21X1_1074 ( .A(_2996_), .B(micro_hash_synth_1_W_13__3_), .C(_2505_), .Y(_2506_) );
	AOI21X1 AOI21X1_757 ( .A(_2996_), .B(micro_hash_synth_1_W_13__3_), .C(_2506_), .Y(_2507_) );
	OAI21X1 OAI21X1_1075 ( .A(_2925__bF_buf4), .B(_2507_), .C(_2504_), .Y(_1436_) );
	NAND2X1 NAND2X1_611 ( .A(micro_hash_synth_1_W_22__4_), .B(_2459__bF_buf0), .Y(_2508_) );
	INVX1 INVX1_897 ( .A(micro_hash_synth_1_W_19__4_), .Y(_2509_) );
	OAI21X1 OAI21X1_1076 ( .A(_2998_), .B(micro_hash_synth_1_W_13__4_), .C(_2509_), .Y(_2510_) );
	AOI21X1 AOI21X1_758 ( .A(_2998_), .B(micro_hash_synth_1_W_13__4_), .C(_2510_), .Y(_2511_) );
	OAI21X1 OAI21X1_1077 ( .A(_2925__bF_buf3), .B(_2511_), .C(_2508_), .Y(_1437_) );
	NAND2X1 NAND2X1_612 ( .A(micro_hash_synth_1_W_22__5_), .B(_2459__bF_buf6), .Y(_2512_) );
	INVX1 INVX1_898 ( .A(micro_hash_synth_1_W_19__5_), .Y(_2513_) );
	OAI21X1 OAI21X1_1078 ( .A(_3000_), .B(micro_hash_synth_1_W_13__5_), .C(_2513_), .Y(_2514_) );
	AOI21X1 AOI21X1_759 ( .A(_3000_), .B(micro_hash_synth_1_W_13__5_), .C(_2514_), .Y(_2515_) );
	OAI21X1 OAI21X1_1079 ( .A(_2925__bF_buf2), .B(_2515_), .C(_2512_), .Y(_1438_) );
	NAND2X1 NAND2X1_613 ( .A(micro_hash_synth_1_W_22__6_), .B(_2459__bF_buf5), .Y(_2516_) );
	INVX1 INVX1_899 ( .A(micro_hash_synth_1_W_19__6_), .Y(_2517_) );
	OAI21X1 OAI21X1_1080 ( .A(_3002_), .B(micro_hash_synth_1_W_13__6_), .C(_2517_), .Y(_2518_) );
	AOI21X1 AOI21X1_760 ( .A(_3002_), .B(micro_hash_synth_1_W_13__6_), .C(_2518_), .Y(_2519_) );
	OAI21X1 OAI21X1_1081 ( .A(_2925__bF_buf1), .B(_2519_), .C(_2516_), .Y(_1439_) );
	NAND2X1 NAND2X1_614 ( .A(micro_hash_synth_1_W_22__7_), .B(_2459__bF_buf4), .Y(_2520_) );
	INVX1 INVX1_900 ( .A(micro_hash_synth_1_W_19__7_), .Y(_2521_) );
	OAI21X1 OAI21X1_1082 ( .A(_3004_), .B(micro_hash_synth_1_W_13__7_), .C(_2521_), .Y(_2522_) );
	AOI21X1 AOI21X1_761 ( .A(_3004_), .B(micro_hash_synth_1_W_13__7_), .C(_2522_), .Y(_2523_) );
	OAI21X1 OAI21X1_1083 ( .A(_2925__bF_buf0), .B(_2523_), .C(_2520_), .Y(_1440_) );
	INVX1 INVX1_901 ( .A(bloque_in_72_), .Y(_2524_) );
	NAND2X1 NAND2X1_615 ( .A(micro_hash_synth_1_W_9__0_), .B(_2459__bF_buf3), .Y(_2525_) );
	OAI21X1 OAI21X1_1084 ( .A(_2524_), .B(_2925__bF_buf15), .C(_2525_), .Y(_1441_) );
	INVX1 INVX1_902 ( .A(bloque_in_73_), .Y(_2526_) );
	NAND2X1 NAND2X1_616 ( .A(micro_hash_synth_1_W_9__1_), .B(_2459__bF_buf2), .Y(_2527_) );
	OAI21X1 OAI21X1_1085 ( .A(_2526_), .B(_2925__bF_buf14), .C(_2527_), .Y(_1442_) );
	INVX1 INVX1_903 ( .A(bloque_in_74_), .Y(_2528_) );
	NAND2X1 NAND2X1_617 ( .A(micro_hash_synth_1_W_9__2_), .B(_2459__bF_buf1), .Y(_2529_) );
	OAI21X1 OAI21X1_1086 ( .A(_2528_), .B(_2925__bF_buf13), .C(_2529_), .Y(_1443_) );
	INVX1 INVX1_904 ( .A(bloque_in_75_), .Y(_2530_) );
	NAND2X1 NAND2X1_618 ( .A(micro_hash_synth_1_W_9__3_), .B(_2459__bF_buf0), .Y(_2531_) );
	OAI21X1 OAI21X1_1087 ( .A(_2530_), .B(_2925__bF_buf12), .C(_2531_), .Y(_1444_) );
	INVX1 INVX1_905 ( .A(bloque_in_76_), .Y(_2532_) );
	NAND2X1 NAND2X1_619 ( .A(micro_hash_synth_1_W_9__4_), .B(_2459__bF_buf6), .Y(_2533_) );
	OAI21X1 OAI21X1_1088 ( .A(_2532_), .B(_2925__bF_buf11), .C(_2533_), .Y(_1446_) );
	INVX1 INVX1_906 ( .A(bloque_in_77_), .Y(_2534_) );
	NAND2X1 NAND2X1_620 ( .A(micro_hash_synth_1_W_9__5_), .B(_2459__bF_buf5), .Y(_2535_) );
	OAI21X1 OAI21X1_1089 ( .A(_2534_), .B(_2925__bF_buf10), .C(_2535_), .Y(_1447_) );
	INVX1 INVX1_907 ( .A(bloque_in_78_), .Y(_2536_) );
	OAI22X1 OAI22X1_331 ( .A(_2536_), .B(_2925__bF_buf9), .C(_2930__bF_buf0), .D(_2202_), .Y(_1448_) );
	INVX1 INVX1_908 ( .A(bloque_in_79_), .Y(_2537_) );
	NAND2X1 NAND2X1_621 ( .A(micro_hash_synth_1_W_9__7_), .B(_2459__bF_buf4), .Y(_2538_) );
	OAI21X1 OAI21X1_1090 ( .A(_2537_), .B(_2925__bF_buf8), .C(_2538_), .Y(_1449_) );
	INVX1 INVX1_909 ( .A(micro_hash_synth_1_W_4__0_), .Y(_2539_) );
	INVX1 INVX1_910 ( .A(bloque_in_32_), .Y(_2540_) );
	OAI22X1 OAI22X1_332 ( .A(_2540_), .B(_2925__bF_buf7), .C(_2930__bF_buf13), .D(_2539_), .Y(_1450_) );
	INVX1 INVX1_911 ( .A(micro_hash_synth_1_W_4__1_), .Y(_2541_) );
	INVX1 INVX1_912 ( .A(bloque_in_33_), .Y(_2542_) );
	OAI22X1 OAI22X1_333 ( .A(_2542_), .B(_2925__bF_buf6), .C(_2930__bF_buf12), .D(_2541_), .Y(_1451_) );
	INVX1 INVX1_913 ( .A(micro_hash_synth_1_W_4__2_), .Y(_2543_) );
	INVX1 INVX1_914 ( .A(bloque_in_34_), .Y(_2544_) );
	OAI22X1 OAI22X1_334 ( .A(_2544_), .B(_2925__bF_buf5), .C(_2930__bF_buf11), .D(_2543_), .Y(_1452_) );
	INVX1 INVX1_915 ( .A(micro_hash_synth_1_W_4__3_), .Y(_2545_) );
	INVX1 INVX1_916 ( .A(bloque_in_35_), .Y(_2546_) );
	OAI22X1 OAI22X1_335 ( .A(_2546_), .B(_2925__bF_buf4), .C(_2930__bF_buf10), .D(_2545_), .Y(_1453_) );
	INVX1 INVX1_917 ( .A(micro_hash_synth_1_W_4__4_), .Y(_2547_) );
	INVX1 INVX1_918 ( .A(bloque_in_36_), .Y(_2548_) );
	OAI22X1 OAI22X1_336 ( .A(_2548_), .B(_2925__bF_buf3), .C(_2930__bF_buf9), .D(_2547_), .Y(_1454_) );
	INVX1 INVX1_919 ( .A(micro_hash_synth_1_W_4__5_), .Y(_2549_) );
	INVX1 INVX1_920 ( .A(bloque_in_37_), .Y(_2550_) );
	OAI22X1 OAI22X1_337 ( .A(_2550_), .B(_2925__bF_buf2), .C(_2930__bF_buf8), .D(_2549_), .Y(_1455_) );
	INVX1 INVX1_921 ( .A(micro_hash_synth_1_W_4__6_), .Y(_2551_) );
	INVX1 INVX1_922 ( .A(bloque_in_38_), .Y(_2552_) );
	OAI22X1 OAI22X1_338 ( .A(_2552_), .B(_2925__bF_buf1), .C(_2930__bF_buf7), .D(_2551_), .Y(_1457_) );
	INVX1 INVX1_923 ( .A(micro_hash_synth_1_W_4__7_), .Y(_2553_) );
	INVX1 INVX1_924 ( .A(bloque_in_39_), .Y(_2554_) );
	OAI22X1 OAI22X1_339 ( .A(_2554_), .B(_2925__bF_buf0), .C(_2930__bF_buf6), .D(_2553_), .Y(_1458_) );
	NAND2X1 NAND2X1_622 ( .A(micro_hash_synth_1_W_21__0_), .B(_2459__bF_buf3), .Y(_2555_) );
	OAI21X1 OAI21X1_1091 ( .A(_2481_), .B(micro_hash_synth_1_W_12__0_), .C(_1670_), .Y(_2556_) );
	AOI21X1 AOI21X1_762 ( .A(micro_hash_synth_1_W_12__0_), .B(_2481_), .C(_2556_), .Y(_2557_) );
	OAI21X1 OAI21X1_1092 ( .A(_2925__bF_buf15), .B(_2557_), .C(_2555_), .Y(_1459_) );
	OAI21X1 OAI21X1_1093 ( .A(_1750_), .B(micro_hash_synth_1_W_12__1_), .C(_1703_), .Y(_2558_) );
	AOI21X1 AOI21X1_763 ( .A(micro_hash_synth_1_W_12__1_), .B(_1750_), .C(_2558_), .Y(_2559_) );
	OAI22X1 OAI22X1_340 ( .A(_2925__bF_buf14), .B(_2559_), .C(_2930__bF_buf5), .D(_2437_), .Y(_1460_) );
	OAI21X1 OAI21X1_1094 ( .A(_1884_), .B(micro_hash_synth_1_W_12__2_), .C(_1804_), .Y(_2560_) );
	AOI21X1 AOI21X1_764 ( .A(micro_hash_synth_1_W_12__2_), .B(_1884_), .C(_2560_), .Y(_2561_) );
	OAI22X1 OAI22X1_341 ( .A(_2925__bF_buf13), .B(_2561_), .C(_2930__bF_buf4), .D(_2440_), .Y(_1461_) );
	OAI21X1 OAI21X1_1095 ( .A(_2485_), .B(micro_hash_synth_1_W_12__3_), .C(_1934_), .Y(_2562_) );
	AOI21X1 AOI21X1_765 ( .A(micro_hash_synth_1_W_12__3_), .B(_2485_), .C(_2562_), .Y(_2563_) );
	OAI22X1 OAI22X1_342 ( .A(_2925__bF_buf12), .B(_2563_), .C(_2930__bF_buf3), .D(_2443_), .Y(_1462_) );
	OAI21X1 OAI21X1_1096 ( .A(_2487_), .B(micro_hash_synth_1_W_12__4_), .C(_2031_), .Y(_2564_) );
	AOI21X1 AOI21X1_766 ( .A(micro_hash_synth_1_W_12__4_), .B(_2487_), .C(_2564_), .Y(_2565_) );
	OAI22X1 OAI22X1_343 ( .A(_2925__bF_buf11), .B(_2565_), .C(_2930__bF_buf2), .D(_2446_), .Y(_1463_) );
	OAI21X1 OAI21X1_1097 ( .A(_2489_), .B(micro_hash_synth_1_W_12__5_), .C(_2088_), .Y(_2566_) );
	AOI21X1 AOI21X1_767 ( .A(micro_hash_synth_1_W_12__5_), .B(_2489_), .C(_2566_), .Y(_2567_) );
	OAI22X1 OAI22X1_344 ( .A(_2925__bF_buf10), .B(_2567_), .C(_2930__bF_buf1), .D(_2449_), .Y(_1464_) );
	OAI21X1 OAI21X1_1098 ( .A(_2212_), .B(micro_hash_synth_1_W_12__6_), .C(_2172_), .Y(_2568_) );
	AOI21X1 AOI21X1_768 ( .A(micro_hash_synth_1_W_12__6_), .B(_2212_), .C(_2568_), .Y(_2569_) );
	OAI22X1 OAI22X1_345 ( .A(_2925__bF_buf9), .B(_2569_), .C(_2930__bF_buf0), .D(_2452_), .Y(_1465_) );
	OAI21X1 OAI21X1_1099 ( .A(_2492_), .B(micro_hash_synth_1_W_12__7_), .C(_2242_), .Y(_2570_) );
	AOI21X1 AOI21X1_769 ( .A(micro_hash_synth_1_W_12__7_), .B(_2492_), .C(_2570_), .Y(_2571_) );
	OAI22X1 OAI22X1_346 ( .A(_2925__bF_buf8), .B(_2571_), .C(_2930__bF_buf13), .D(_2456_), .Y(_1466_) );
	NAND2X1 NAND2X1_623 ( .A(micro_hash_synth_1_W_20__0_), .B(_2459__bF_buf2), .Y(_2572_) );
	INVX1 INVX1_925 ( .A(micro_hash_synth_1_W_6__0_), .Y(_2573_) );
	INVX1 INVX1_926 ( .A(micro_hash_synth_1_W_17__0_), .Y(_2574_) );
	OAI21X1 OAI21X1_1100 ( .A(_2573_), .B(micro_hash_synth_1_W_11__0_), .C(_2574_), .Y(_2575_) );
	AOI21X1 AOI21X1_770 ( .A(micro_hash_synth_1_W_11__0_), .B(_2573_), .C(_2575_), .Y(_2576_) );
	OAI21X1 OAI21X1_1101 ( .A(_2925__bF_buf7), .B(_2576_), .C(_2572_), .Y(_1468_) );
	NAND2X1 NAND2X1_624 ( .A(micro_hash_synth_1_W_20__1_), .B(_2459__bF_buf1), .Y(_2577_) );
	INVX1 INVX1_927 ( .A(micro_hash_synth_1_W_6__1_), .Y(_2578_) );
	INVX1 INVX1_928 ( .A(micro_hash_synth_1_W_17__1_), .Y(_2579_) );
	OAI21X1 OAI21X1_1102 ( .A(_2578_), .B(micro_hash_synth_1_W_11__1_), .C(_2579_), .Y(_2580_) );
	AOI21X1 AOI21X1_771 ( .A(micro_hash_synth_1_W_11__1_), .B(_2578_), .C(_2580_), .Y(_2581_) );
	OAI21X1 OAI21X1_1103 ( .A(_2925__bF_buf6), .B(_2581_), .C(_2577_), .Y(_1469_) );
	NAND2X1 NAND2X1_625 ( .A(micro_hash_synth_1_W_20__2_), .B(_2459__bF_buf0), .Y(_2582_) );
	INVX1 INVX1_929 ( .A(micro_hash_synth_1_W_6__2_), .Y(_2583_) );
	INVX1 INVX1_930 ( .A(micro_hash_synth_1_W_17__2_), .Y(_2584_) );
	OAI21X1 OAI21X1_1104 ( .A(_2583_), .B(micro_hash_synth_1_W_11__2_), .C(_2584_), .Y(_2585_) );
	AOI21X1 AOI21X1_772 ( .A(micro_hash_synth_1_W_11__2_), .B(_2583_), .C(_2585_), .Y(_2586_) );
	OAI21X1 OAI21X1_1105 ( .A(_2925__bF_buf5), .B(_2586_), .C(_2582_), .Y(_1470_) );
	NAND2X1 NAND2X1_626 ( .A(micro_hash_synth_1_W_20__3_), .B(_2459__bF_buf6), .Y(_2587_) );
	INVX1 INVX1_931 ( .A(micro_hash_synth_1_W_6__3_), .Y(_2588_) );
	INVX1 INVX1_932 ( .A(micro_hash_synth_1_W_17__3_), .Y(_2589_) );
	OAI21X1 OAI21X1_1106 ( .A(_2588_), .B(micro_hash_synth_1_W_11__3_), .C(_2589_), .Y(_2590_) );
	AOI21X1 AOI21X1_773 ( .A(micro_hash_synth_1_W_11__3_), .B(_2588_), .C(_2590_), .Y(_2591_) );
	OAI21X1 OAI21X1_1107 ( .A(_2925__bF_buf4), .B(_2591_), .C(_2587_), .Y(_1471_) );
	NAND2X1 NAND2X1_627 ( .A(micro_hash_synth_1_W_20__4_), .B(_2459__bF_buf5), .Y(_2592_) );
	INVX1 INVX1_933 ( .A(micro_hash_synth_1_W_6__4_), .Y(_2593_) );
	INVX1 INVX1_934 ( .A(micro_hash_synth_1_W_17__4_), .Y(_2594_) );
	OAI21X1 OAI21X1_1108 ( .A(_2593_), .B(micro_hash_synth_1_W_11__4_), .C(_2594_), .Y(_2595_) );
	AOI21X1 AOI21X1_774 ( .A(micro_hash_synth_1_W_11__4_), .B(_2593_), .C(_2595_), .Y(_2596_) );
	OAI21X1 OAI21X1_1109 ( .A(_2925__bF_buf3), .B(_2596_), .C(_2592_), .Y(_1472_) );
	NAND2X1 NAND2X1_628 ( .A(micro_hash_synth_1_W_20__5_), .B(_2459__bF_buf4), .Y(_2597_) );
	INVX1 INVX1_935 ( .A(micro_hash_synth_1_W_6__5_), .Y(_2598_) );
	INVX1 INVX1_936 ( .A(micro_hash_synth_1_W_17__5_), .Y(_2599_) );
	OAI21X1 OAI21X1_1110 ( .A(_2598_), .B(micro_hash_synth_1_W_11__5_), .C(_2599_), .Y(_2600_) );
	AOI21X1 AOI21X1_775 ( .A(micro_hash_synth_1_W_11__5_), .B(_2598_), .C(_2600_), .Y(_2601_) );
	OAI21X1 OAI21X1_1111 ( .A(_2925__bF_buf2), .B(_2601_), .C(_2597_), .Y(_1473_) );
	INVX1 INVX1_937 ( .A(micro_hash_synth_1_W_6__6_), .Y(_2602_) );
	INVX1 INVX1_938 ( .A(micro_hash_synth_1_W_17__6_), .Y(_2603_) );
	OAI21X1 OAI21X1_1112 ( .A(_2602_), .B(micro_hash_synth_1_W_11__6_), .C(_2603_), .Y(_2604_) );
	AOI21X1 AOI21X1_776 ( .A(micro_hash_synth_1_W_11__6_), .B(_2602_), .C(_2604_), .Y(_2605_) );
	OAI22X1 OAI22X1_347 ( .A(_2925__bF_buf1), .B(_2605_), .C(_2930__bF_buf12), .D(_2476_), .Y(_1474_) );
	NAND2X1 NAND2X1_629 ( .A(micro_hash_synth_1_W_20__7_), .B(_2459__bF_buf3), .Y(_2606_) );
	INVX1 INVX1_939 ( .A(micro_hash_synth_1_W_17__7_), .Y(_2607_) );
	OAI21X1 OAI21X1_1113 ( .A(_2280_), .B(micro_hash_synth_1_W_11__7_), .C(_2607_), .Y(_2608_) );
	AOI21X1 AOI21X1_777 ( .A(micro_hash_synth_1_W_11__7_), .B(_2280_), .C(_2608_), .Y(_2609_) );
	OAI21X1 OAI21X1_1114 ( .A(_2925__bF_buf0), .B(_2609_), .C(_2606_), .Y(_1475_) );
	INVX1 INVX1_940 ( .A(bloque_in_96_), .Y(_2610_) );
	NAND2X1 NAND2X1_630 ( .A(micro_hash_synth_1_W_12__0_), .B(_2459__bF_buf2), .Y(_2611_) );
	OAI21X1 OAI21X1_1115 ( .A(_2610_), .B(_2925__bF_buf15), .C(_2611_), .Y(_1476_) );
	INVX1 INVX1_941 ( .A(bloque_in_97_), .Y(_2612_) );
	OAI22X1 OAI22X1_348 ( .A(_2612_), .B(_2925__bF_buf14), .C(_2930__bF_buf11), .D(_2934_), .Y(_1477_) );
	INVX1 INVX1_942 ( .A(bloque_in_98_), .Y(_2613_) );
	OAI22X1 OAI22X1_349 ( .A(_2613_), .B(_2925__bF_buf13), .C(_2930__bF_buf10), .D(_2939_), .Y(_1479_) );
	INVX1 INVX1_943 ( .A(bloque_in_99_), .Y(_2614_) );
	NAND2X1 NAND2X1_631 ( .A(micro_hash_synth_1_W_12__3_), .B(_2459__bF_buf1), .Y(_2615_) );
	OAI21X1 OAI21X1_1116 ( .A(_2614_), .B(_2925__bF_buf12), .C(_2615_), .Y(_1480_) );
	INVX1 INVX1_944 ( .A(bloque_in_100_), .Y(_2616_) );
	NAND2X1 NAND2X1_632 ( .A(micro_hash_synth_1_W_12__4_), .B(_2459__bF_buf0), .Y(_2617_) );
	OAI21X1 OAI21X1_1117 ( .A(_2616_), .B(_2925__bF_buf11), .C(_2617_), .Y(_1481_) );
	INVX1 INVX1_945 ( .A(bloque_in_101_), .Y(_2618_) );
	NAND2X1 NAND2X1_633 ( .A(micro_hash_synth_1_W_12__5_), .B(_2459__bF_buf6), .Y(_2619_) );
	OAI21X1 OAI21X1_1118 ( .A(_2618_), .B(_2925__bF_buf10), .C(_2619_), .Y(_1482_) );
	INVX1 INVX1_946 ( .A(bloque_in_102_), .Y(_2620_) );
	OAI22X1 OAI22X1_350 ( .A(_2620_), .B(_2925__bF_buf9), .C(_2930__bF_buf9), .D(_2953_), .Y(_1483_) );
	INVX1 INVX1_947 ( .A(bloque_in_103_), .Y(_2621_) );
	OAI22X1 OAI22X1_351 ( .A(_2621_), .B(_2925__bF_buf8), .C(_2930__bF_buf8), .D(_2958_), .Y(_1484_) );
	INVX1 INVX1_948 ( .A(micro_hash_synth_1_W_5__0_), .Y(_2622_) );
	OAI21X1 OAI21X1_1119 ( .A(_2622_), .B(micro_hash_synth_1_W_10__0_), .C(_1673_), .Y(_2623_) );
	AOI21X1 AOI21X1_778 ( .A(_2622_), .B(micro_hash_synth_1_W_10__0_), .C(_2623_), .Y(_2624_) );
	OAI22X1 OAI22X1_352 ( .A(_2925__bF_buf7), .B(_2624_), .C(_2930__bF_buf7), .D(_2495_), .Y(_1488_) );
	OAI21X1 OAI21X1_1120 ( .A(_1745_), .B(micro_hash_synth_1_W_10__1_), .C(_1707_), .Y(_2625_) );
	AOI21X1 AOI21X1_779 ( .A(_1745_), .B(micro_hash_synth_1_W_10__1_), .C(_2625_), .Y(_2626_) );
	OAI22X1 OAI22X1_353 ( .A(_2925__bF_buf6), .B(_2626_), .C(_2930__bF_buf6), .D(_2498_), .Y(_1489_) );
	OAI21X1 OAI21X1_1121 ( .A(_1879_), .B(micro_hash_synth_1_W_10__2_), .C(_1808_), .Y(_2627_) );
	AOI21X1 AOI21X1_780 ( .A(_1879_), .B(micro_hash_synth_1_W_10__2_), .C(_2627_), .Y(_2628_) );
	OAI22X1 OAI22X1_354 ( .A(_2925__bF_buf5), .B(_2628_), .C(_2930__bF_buf5), .D(_2501_), .Y(_1490_) );
	INVX1 INVX1_949 ( .A(micro_hash_synth_1_W_5__3_), .Y(_2629_) );
	OAI21X1 OAI21X1_1122 ( .A(_2629_), .B(micro_hash_synth_1_W_10__3_), .C(_1938_), .Y(_2630_) );
	AOI21X1 AOI21X1_781 ( .A(_2629_), .B(micro_hash_synth_1_W_10__3_), .C(_2630_), .Y(_2631_) );
	OAI22X1 OAI22X1_355 ( .A(_2925__bF_buf4), .B(_2631_), .C(_2930__bF_buf4), .D(_2505_), .Y(_1491_) );
	INVX1 INVX1_950 ( .A(micro_hash_synth_1_W_5__4_), .Y(_2632_) );
	OAI21X1 OAI21X1_1123 ( .A(_2632_), .B(micro_hash_synth_1_W_10__4_), .C(_2035_), .Y(_2633_) );
	AOI21X1 AOI21X1_782 ( .A(_2632_), .B(micro_hash_synth_1_W_10__4_), .C(_2633_), .Y(_2634_) );
	OAI22X1 OAI22X1_356 ( .A(_2925__bF_buf3), .B(_2634_), .C(_2930__bF_buf3), .D(_2509_), .Y(_1493_) );
	INVX1 INVX1_951 ( .A(micro_hash_synth_1_W_5__5_), .Y(_2635_) );
	OAI21X1 OAI21X1_1124 ( .A(_2635_), .B(micro_hash_synth_1_W_10__5_), .C(_2092_), .Y(_2636_) );
	AOI21X1 AOI21X1_783 ( .A(_2635_), .B(micro_hash_synth_1_W_10__5_), .C(_2636_), .Y(_2637_) );
	OAI22X1 OAI22X1_357 ( .A(_2925__bF_buf2), .B(_2637_), .C(_2930__bF_buf2), .D(_2513_), .Y(_1494_) );
	INVX1 INVX1_952 ( .A(micro_hash_synth_1_W_5__6_), .Y(_2638_) );
	OAI21X1 OAI21X1_1125 ( .A(_2638_), .B(micro_hash_synth_1_W_10__6_), .C(_2175_), .Y(_2639_) );
	AOI21X1 AOI21X1_784 ( .A(_2638_), .B(micro_hash_synth_1_W_10__6_), .C(_2639_), .Y(_2640_) );
	OAI22X1 OAI22X1_358 ( .A(_2925__bF_buf1), .B(_2640_), .C(_2930__bF_buf1), .D(_2517_), .Y(_1495_) );
	INVX1 INVX1_953 ( .A(micro_hash_synth_1_W_5__7_), .Y(_2641_) );
	INVX1 INVX1_954 ( .A(micro_hash_synth_1_W_16__7_), .Y(_2642_) );
	OAI21X1 OAI21X1_1126 ( .A(_2641_), .B(micro_hash_synth_1_W_10__7_), .C(_2642_), .Y(_2643_) );
	AOI21X1 AOI21X1_785 ( .A(_2641_), .B(micro_hash_synth_1_W_10__7_), .C(_2643_), .Y(_2644_) );
	OAI22X1 OAI22X1_359 ( .A(_2925__bF_buf0), .B(_2644_), .C(_2930__bF_buf0), .D(_2521_), .Y(_1496_) );
	INVX1 INVX1_955 ( .A(bloque_in_40_), .Y(_2645_) );
	OAI22X1 OAI22X1_360 ( .A(_2645_), .B(_2925__bF_buf15), .C(_2930__bF_buf13), .D(_2622_), .Y(_1246_) );
	INVX1 INVX1_956 ( .A(bloque_in_41_), .Y(_2646_) );
	OAI22X1 OAI22X1_361 ( .A(_2646_), .B(_2925__bF_buf14), .C(_2930__bF_buf12), .D(_1745_), .Y(_1247_) );
	INVX1 INVX1_957 ( .A(bloque_in_42_), .Y(_2647_) );
	OAI22X1 OAI22X1_362 ( .A(_2647_), .B(_2925__bF_buf13), .C(_2930__bF_buf11), .D(_1879_), .Y(_1248_) );
	INVX1 INVX1_958 ( .A(bloque_in_43_), .Y(_2648_) );
	OAI22X1 OAI22X1_363 ( .A(_2648_), .B(_2925__bF_buf12), .C(_2930__bF_buf10), .D(_2629_), .Y(_1249_) );
	INVX1 INVX1_959 ( .A(bloque_in_44_), .Y(_2649_) );
	OAI22X1 OAI22X1_364 ( .A(_2649_), .B(_2925__bF_buf11), .C(_2930__bF_buf9), .D(_2632_), .Y(_1250_) );
	INVX1 INVX1_960 ( .A(bloque_in_45_), .Y(_2650_) );
	OAI22X1 OAI22X1_365 ( .A(_2650_), .B(_2925__bF_buf10), .C(_2930__bF_buf8), .D(_2635_), .Y(_1251_) );
	INVX1 INVX1_961 ( .A(bloque_in_46_), .Y(_2651_) );
	OAI22X1 OAI22X1_366 ( .A(_2651_), .B(_2925__bF_buf9), .C(_2930__bF_buf7), .D(_2638_), .Y(_1252_) );
	INVX1 INVX1_962 ( .A(bloque_in_47_), .Y(_2652_) );
	OAI22X1 OAI22X1_367 ( .A(_2652_), .B(_2925__bF_buf8), .C(_2930__bF_buf6), .D(_2641_), .Y(_1254_) );
	INVX1 INVX1_963 ( .A(micro_hash_synth_1_W_14__0_), .Y(_2653_) );
	INVX1 INVX1_964 ( .A(bloque_in_112_), .Y(_2654_) );
	OAI22X1 OAI22X1_368 ( .A(_2654_), .B(_2925__bF_buf7), .C(_2930__bF_buf5), .D(_2653_), .Y(_1258_) );
	INVX1 INVX1_965 ( .A(micro_hash_synth_1_W_14__1_), .Y(_2655_) );
	INVX1 INVX1_966 ( .A(bloque_in_113_), .Y(_2656_) );
	OAI22X1 OAI22X1_369 ( .A(_2656_), .B(_2925__bF_buf6), .C(_2930__bF_buf4), .D(_2655_), .Y(_1259_) );
	INVX1 INVX1_967 ( .A(micro_hash_synth_1_W_14__2_), .Y(_2657_) );
	INVX1 INVX1_968 ( .A(bloque_in_114_), .Y(_2658_) );
	OAI22X1 OAI22X1_370 ( .A(_2658_), .B(_2925__bF_buf5), .C(_2930__bF_buf3), .D(_2657_), .Y(_1260_) );
	INVX1 INVX1_969 ( .A(micro_hash_synth_1_W_14__3_), .Y(_2659_) );
	INVX1 INVX1_970 ( .A(bloque_in_115_), .Y(_2660_) );
	OAI22X1 OAI22X1_371 ( .A(_2660_), .B(_2925__bF_buf4), .C(_2930__bF_buf2), .D(_2659_), .Y(_1261_) );
	INVX1 INVX1_971 ( .A(micro_hash_synth_1_W_14__4_), .Y(_2661_) );
	INVX1 INVX1_972 ( .A(bloque_in_116_), .Y(_2662_) );
	OAI22X1 OAI22X1_372 ( .A(_2662_), .B(_2925__bF_buf3), .C(_2930__bF_buf1), .D(_2661_), .Y(_1262_) );
	INVX1 INVX1_973 ( .A(micro_hash_synth_1_W_14__5_), .Y(_2663_) );
	INVX1 INVX1_974 ( .A(bloque_in_117_), .Y(_2664_) );
	OAI22X1 OAI22X1_373 ( .A(_2664_), .B(_2925__bF_buf2), .C(_2930__bF_buf0), .D(_2663_), .Y(_1263_) );
	INVX1 INVX1_975 ( .A(micro_hash_synth_1_W_14__6_), .Y(_2665_) );
	INVX1 INVX1_976 ( .A(bloque_in_118_), .Y(_2666_) );
	OAI22X1 OAI22X1_374 ( .A(_2666_), .B(_2925__bF_buf1), .C(_2930__bF_buf13), .D(_2665_), .Y(_1264_) );
	INVX1 INVX1_977 ( .A(micro_hash_synth_1_W_14__7_), .Y(_2667_) );
	INVX1 INVX1_978 ( .A(bloque_in_119_), .Y(_2668_) );
	OAI22X1 OAI22X1_375 ( .A(_2668_), .B(_2925__bF_buf0), .C(_2930__bF_buf12), .D(_2667_), .Y(_1265_) );
	INVX1 INVX1_979 ( .A(bloque_in_0_), .Y(_2669_) );
	OAI22X1 OAI22X1_376 ( .A(_2669_), .B(_2925__bF_buf15), .C(_2930__bF_buf11), .D(_3031_), .Y(_1267_) );
	INVX1 INVX1_980 ( .A(bloque_in_1_), .Y(_2670_) );
	OAI22X1 OAI22X1_377 ( .A(_2670_), .B(_2925__bF_buf14), .C(_2930__bF_buf10), .D(_3032_), .Y(_1268_) );
	INVX1 INVX1_981 ( .A(bloque_in_2_), .Y(_2671_) );
	OAI22X1 OAI22X1_378 ( .A(_2671_), .B(_2925__bF_buf13), .C(_2930__bF_buf9), .D(_3033_), .Y(_1270_) );
	INVX1 INVX1_982 ( .A(bloque_in_3_), .Y(_2672_) );
	OAI22X1 OAI22X1_379 ( .A(_2672_), .B(_2925__bF_buf12), .C(_2930__bF_buf8), .D(_3034_), .Y(_1271_) );
	INVX1 INVX1_983 ( .A(bloque_in_4_), .Y(_2673_) );
	OAI22X1 OAI22X1_380 ( .A(_2673_), .B(_2925__bF_buf11), .C(_2930__bF_buf7), .D(_3035_), .Y(_1272_) );
	INVX1 INVX1_984 ( .A(bloque_in_5_), .Y(_2674_) );
	OAI22X1 OAI22X1_381 ( .A(_2674_), .B(_2925__bF_buf10), .C(_2930__bF_buf6), .D(_3036_), .Y(_1273_) );
	INVX1 INVX1_985 ( .A(bloque_in_6_), .Y(_2675_) );
	OAI22X1 OAI22X1_382 ( .A(_2675_), .B(_2925__bF_buf9), .C(_2930__bF_buf5), .D(_3037_), .Y(_1274_) );
	INVX1 INVX1_986 ( .A(bloque_in_7_), .Y(_2676_) );
	OAI22X1 OAI22X1_383 ( .A(_2676_), .B(_2925__bF_buf8), .C(_2930__bF_buf4), .D(_3038_), .Y(_1275_) );
	INVX1 INVX1_987 ( .A(micro_hash_synth_1_W_15__0_), .Y(_2677_) );
	OAI21X1 OAI21X1_1127 ( .A(_2539_), .B(micro_hash_synth_1_W_9__0_), .C(_2677_), .Y(_2678_) );
	AOI21X1 AOI21X1_786 ( .A(_2539_), .B(micro_hash_synth_1_W_9__0_), .C(_2678_), .Y(_2679_) );
	OAI22X1 OAI22X1_384 ( .A(_2925__bF_buf7), .B(_2679_), .C(_2930__bF_buf3), .D(_1670_), .Y(_1276_) );
	INVX1 INVX1_988 ( .A(micro_hash_synth_1_W_15__1_), .Y(_2680_) );
	OAI21X1 OAI21X1_1128 ( .A(_2541_), .B(micro_hash_synth_1_W_9__1_), .C(_2680_), .Y(_2681_) );
	AOI21X1 AOI21X1_787 ( .A(_2541_), .B(micro_hash_synth_1_W_9__1_), .C(_2681_), .Y(_2682_) );
	OAI22X1 OAI22X1_385 ( .A(_2925__bF_buf6), .B(_2682_), .C(_2930__bF_buf2), .D(_1703_), .Y(_1277_) );
	INVX1 INVX1_989 ( .A(micro_hash_synth_1_W_15__2_), .Y(_2683_) );
	OAI21X1 OAI21X1_1129 ( .A(_2543_), .B(micro_hash_synth_1_W_9__2_), .C(_2683_), .Y(_2684_) );
	AOI21X1 AOI21X1_788 ( .A(_2543_), .B(micro_hash_synth_1_W_9__2_), .C(_2684_), .Y(_2685_) );
	OAI22X1 OAI22X1_386 ( .A(_2925__bF_buf5), .B(_2685_), .C(_2930__bF_buf1), .D(_1804_), .Y(_1278_) );
	INVX1 INVX1_990 ( .A(micro_hash_synth_1_W_15__3_), .Y(_2686_) );
	OAI21X1 OAI21X1_1130 ( .A(_2545_), .B(micro_hash_synth_1_W_9__3_), .C(_2686_), .Y(_2687_) );
	AOI21X1 AOI21X1_789 ( .A(_2545_), .B(micro_hash_synth_1_W_9__3_), .C(_2687_), .Y(_2688_) );
	OAI22X1 OAI22X1_387 ( .A(_2925__bF_buf4), .B(_2688_), .C(_2930__bF_buf0), .D(_1934_), .Y(_1279_) );
	INVX1 INVX1_991 ( .A(micro_hash_synth_1_W_15__4_), .Y(_2689_) );
	OAI21X1 OAI21X1_1131 ( .A(_2547_), .B(micro_hash_synth_1_W_9__4_), .C(_2689_), .Y(_2690_) );
	AOI21X1 AOI21X1_790 ( .A(_2547_), .B(micro_hash_synth_1_W_9__4_), .C(_2690_), .Y(_2691_) );
	OAI22X1 OAI22X1_388 ( .A(_2925__bF_buf3), .B(_2691_), .C(_2930__bF_buf13), .D(_2031_), .Y(_1280_) );
	INVX1 INVX1_992 ( .A(micro_hash_synth_1_W_15__5_), .Y(_2692_) );
	OAI21X1 OAI21X1_1132 ( .A(_2549_), .B(micro_hash_synth_1_W_9__5_), .C(_2692_), .Y(_2693_) );
	AOI21X1 AOI21X1_791 ( .A(_2549_), .B(micro_hash_synth_1_W_9__5_), .C(_2693_), .Y(_2694_) );
	OAI22X1 OAI22X1_389 ( .A(_2925__bF_buf2), .B(_2694_), .C(_2930__bF_buf12), .D(_2088_), .Y(_1281_) );
	OAI21X1 OAI21X1_1133 ( .A(_2551_), .B(micro_hash_synth_1_W_9__6_), .C(_2197_), .Y(_2695_) );
	AOI21X1 AOI21X1_792 ( .A(_2551_), .B(micro_hash_synth_1_W_9__6_), .C(_2695_), .Y(_2696_) );
	OAI22X1 OAI22X1_390 ( .A(_2925__bF_buf1), .B(_2696_), .C(_2930__bF_buf11), .D(_2172_), .Y(_1282_) );
	OAI21X1 OAI21X1_1134 ( .A(_2553_), .B(micro_hash_synth_1_W_9__7_), .C(_2266_), .Y(_2697_) );
	AOI21X1 AOI21X1_793 ( .A(_2553_), .B(micro_hash_synth_1_W_9__7_), .C(_2697_), .Y(_2698_) );
	OAI22X1 OAI22X1_391 ( .A(_2925__bF_buf0), .B(_2698_), .C(_2930__bF_buf10), .D(_2242_), .Y(_1283_) );
	OAI21X1 OAI21X1_1135 ( .A(_3006_), .B(micro_hash_synth_1_W_8__0_), .C(_2653_), .Y(_2699_) );
	AOI21X1 AOI21X1_794 ( .A(micro_hash_synth_1_W_8__0_), .B(_3006_), .C(_2699_), .Y(_2700_) );
	OAI22X1 OAI22X1_392 ( .A(_2925__bF_buf15), .B(_2700_), .C(_2930__bF_buf9), .D(_2574_), .Y(_1284_) );
	OAI21X1 OAI21X1_1136 ( .A(_3008_), .B(micro_hash_synth_1_W_8__1_), .C(_2655_), .Y(_2701_) );
	AOI21X1 AOI21X1_795 ( .A(micro_hash_synth_1_W_8__1_), .B(_3008_), .C(_2701_), .Y(_2702_) );
	OAI22X1 OAI22X1_393 ( .A(_2925__bF_buf14), .B(_2702_), .C(_2930__bF_buf8), .D(_2579_), .Y(_1286_) );
	OAI21X1 OAI21X1_1137 ( .A(_3010_), .B(micro_hash_synth_1_W_8__2_), .C(_2657_), .Y(_2703_) );
	AOI21X1 AOI21X1_796 ( .A(micro_hash_synth_1_W_8__2_), .B(_3010_), .C(_2703_), .Y(_2704_) );
	OAI22X1 OAI22X1_394 ( .A(_2925__bF_buf13), .B(_2704_), .C(_2930__bF_buf7), .D(_2584_), .Y(_1287_) );
	OAI21X1 OAI21X1_1138 ( .A(_3012_), .B(micro_hash_synth_1_W_8__3_), .C(_2659_), .Y(_2705_) );
	AOI21X1 AOI21X1_797 ( .A(micro_hash_synth_1_W_8__3_), .B(_3012_), .C(_2705_), .Y(_2706_) );
	OAI22X1 OAI22X1_395 ( .A(_2925__bF_buf12), .B(_2706_), .C(_2930__bF_buf6), .D(_2589_), .Y(_1288_) );
	OAI21X1 OAI21X1_1139 ( .A(_3014_), .B(micro_hash_synth_1_W_8__4_), .C(_2661_), .Y(_2707_) );
	AOI21X1 AOI21X1_798 ( .A(micro_hash_synth_1_W_8__4_), .B(_3014_), .C(_2707_), .Y(_2708_) );
	OAI22X1 OAI22X1_396 ( .A(_2925__bF_buf11), .B(_2708_), .C(_2930__bF_buf5), .D(_2594_), .Y(_1289_) );
	OAI21X1 OAI21X1_1140 ( .A(_3016_), .B(micro_hash_synth_1_W_8__5_), .C(_2663_), .Y(_2709_) );
	AOI21X1 AOI21X1_799 ( .A(micro_hash_synth_1_W_8__5_), .B(_3016_), .C(_2709_), .Y(_2710_) );
	OAI22X1 OAI22X1_397 ( .A(_2925__bF_buf10), .B(_2710_), .C(_2930__bF_buf4), .D(_2599_), .Y(_1290_) );
	OAI21X1 OAI21X1_1141 ( .A(_3018_), .B(micro_hash_synth_1_W_8__6_), .C(_2665_), .Y(_2711_) );
	AOI21X1 AOI21X1_800 ( .A(micro_hash_synth_1_W_8__6_), .B(_3018_), .C(_2711_), .Y(_2712_) );
	OAI22X1 OAI22X1_398 ( .A(_2925__bF_buf9), .B(_2712_), .C(_2930__bF_buf3), .D(_2603_), .Y(_1291_) );
	OAI21X1 OAI21X1_1142 ( .A(_3020_), .B(micro_hash_synth_1_W_8__7_), .C(_2667_), .Y(_2713_) );
	AOI21X1 AOI21X1_801 ( .A(micro_hash_synth_1_W_8__7_), .B(_3020_), .C(_2713_), .Y(_2714_) );
	OAI22X1 OAI22X1_399 ( .A(_2925__bF_buf8), .B(_2714_), .C(_2930__bF_buf2), .D(_2607_), .Y(_1292_) );
	INVX1 INVX1_993 ( .A(bloque_in_120_), .Y(_2715_) );
	OAI22X1 OAI22X1_400 ( .A(_2715_), .B(_2925__bF_buf7), .C(_2930__bF_buf1), .D(_2677_), .Y(_1293_) );
	INVX1 INVX1_994 ( .A(bloque_in_121_), .Y(_2716_) );
	OAI22X1 OAI22X1_401 ( .A(_2716_), .B(_2925__bF_buf6), .C(_2930__bF_buf0), .D(_2680_), .Y(_1294_) );
	INVX1 INVX1_995 ( .A(bloque_in_122_), .Y(_2717_) );
	OAI22X1 OAI22X1_402 ( .A(_2717_), .B(_2925__bF_buf5), .C(_2930__bF_buf13), .D(_2683_), .Y(_1295_) );
	INVX1 INVX1_996 ( .A(bloque_in_123_), .Y(_2718_) );
	OAI22X1 OAI22X1_403 ( .A(_2718_), .B(_2925__bF_buf4), .C(_2930__bF_buf12), .D(_2686_), .Y(_1296_) );
	INVX1 INVX1_997 ( .A(bloque_in_124_), .Y(_2719_) );
	OAI22X1 OAI22X1_404 ( .A(_2719_), .B(_2925__bF_buf3), .C(_2930__bF_buf11), .D(_2689_), .Y(_1297_) );
	INVX1 INVX1_998 ( .A(bloque_in_125_), .Y(_2720_) );
	OAI22X1 OAI22X1_405 ( .A(_2720_), .B(_2925__bF_buf2), .C(_2930__bF_buf10), .D(_2692_), .Y(_1298_) );
	INVX1 INVX1_999 ( .A(bloque_in_126_), .Y(_2721_) );
	OAI22X1 OAI22X1_406 ( .A(_2721_), .B(_2925__bF_buf1), .C(_2930__bF_buf9), .D(_2197_), .Y(_1299_) );
	INVX1 INVX1_1000 ( .A(bloque_in_127_), .Y(_2722_) );
	OAI22X1 OAI22X1_407 ( .A(_2722_), .B(_2925__bF_buf0), .C(_2930__bF_buf8), .D(_2266_), .Y(_1300_) );
	INVX1 INVX1_1001 ( .A(bloque_in_48_), .Y(_2723_) );
	OAI22X1 OAI22X1_408 ( .A(_2723_), .B(_2925__bF_buf15), .C(_2930__bF_buf7), .D(_2573_), .Y(_1302_) );
	INVX1 INVX1_1002 ( .A(bloque_in_49_), .Y(_2724_) );
	OAI22X1 OAI22X1_409 ( .A(_2724_), .B(_2925__bF_buf14), .C(_2930__bF_buf6), .D(_2578_), .Y(_1303_) );
	INVX1 INVX1_1003 ( .A(bloque_in_50_), .Y(_2725_) );
	OAI22X1 OAI22X1_410 ( .A(_2725_), .B(_2925__bF_buf13), .C(_2930__bF_buf5), .D(_2583_), .Y(_1304_) );
	INVX1 INVX1_1004 ( .A(bloque_in_51_), .Y(_2726_) );
	OAI22X1 OAI22X1_411 ( .A(_2726_), .B(_2925__bF_buf12), .C(_2930__bF_buf4), .D(_2588_), .Y(_1305_) );
	INVX1 INVX1_1005 ( .A(bloque_in_52_), .Y(_2727_) );
	OAI22X1 OAI22X1_412 ( .A(_2727_), .B(_2925__bF_buf11), .C(_2930__bF_buf3), .D(_2593_), .Y(_1306_) );
	INVX1 INVX1_1006 ( .A(bloque_in_53_), .Y(_2728_) );
	OAI22X1 OAI22X1_413 ( .A(_2728_), .B(_2925__bF_buf10), .C(_2930__bF_buf2), .D(_2598_), .Y(_1307_) );
	INVX1 INVX1_1007 ( .A(bloque_in_54_), .Y(_2729_) );
	OAI22X1 OAI22X1_414 ( .A(_2729_), .B(_2925__bF_buf9), .C(_2930__bF_buf1), .D(_2602_), .Y(_1308_) );
	INVX1 INVX1_1008 ( .A(bloque_in_55_), .Y(_2730_) );
	OAI22X1 OAI22X1_415 ( .A(_2730_), .B(_2925__bF_buf8), .C(_2930__bF_buf0), .D(_2280_), .Y(_1309_) );
	INVX1 INVX1_1009 ( .A(micro_hash_synth_1_W_13__0_), .Y(_2731_) );
	INVX1 INVX1_1010 ( .A(bloque_in_104_), .Y(_2732_) );
	OAI22X1 OAI22X1_416 ( .A(_2732_), .B(_2925__bF_buf7), .C(_2930__bF_buf13), .D(_2731_), .Y(_1310_) );
	INVX1 INVX1_1011 ( .A(micro_hash_synth_1_W_13__1_), .Y(_2733_) );
	INVX1 INVX1_1012 ( .A(bloque_in_105_), .Y(_2734_) );
	OAI22X1 OAI22X1_417 ( .A(_2734_), .B(_2925__bF_buf6), .C(_2930__bF_buf12), .D(_2733_), .Y(_1311_) );
	INVX1 INVX1_1013 ( .A(micro_hash_synth_1_W_13__2_), .Y(_2735_) );
	INVX1 INVX1_1014 ( .A(bloque_in_106_), .Y(_2736_) );
	OAI22X1 OAI22X1_418 ( .A(_2736_), .B(_2925__bF_buf5), .C(_2930__bF_buf11), .D(_2735_), .Y(_1312_) );
	INVX1 INVX1_1015 ( .A(micro_hash_synth_1_W_13__3_), .Y(_2737_) );
	INVX1 INVX1_1016 ( .A(bloque_in_107_), .Y(_2738_) );
	OAI22X1 OAI22X1_419 ( .A(_2738_), .B(_2925__bF_buf4), .C(_2930__bF_buf10), .D(_2737_), .Y(_1313_) );
	INVX1 INVX1_1017 ( .A(micro_hash_synth_1_W_13__4_), .Y(_2739_) );
	INVX1 INVX1_1018 ( .A(bloque_in_108_), .Y(_2740_) );
	OAI22X1 OAI22X1_420 ( .A(_2740_), .B(_2925__bF_buf3), .C(_2930__bF_buf9), .D(_2739_), .Y(_1314_) );
	INVX1 INVX1_1019 ( .A(micro_hash_synth_1_W_13__5_), .Y(_2741_) );
	INVX1 INVX1_1020 ( .A(bloque_in_109_), .Y(_2742_) );
	OAI22X1 OAI22X1_421 ( .A(_2742_), .B(_2925__bF_buf2), .C(_2930__bF_buf8), .D(_2741_), .Y(_1315_) );
	INVX1 INVX1_1021 ( .A(micro_hash_synth_1_W_13__6_), .Y(_2743_) );
	INVX1 INVX1_1022 ( .A(bloque_in_110_), .Y(_2744_) );
	OAI22X1 OAI22X1_422 ( .A(_2744_), .B(_2925__bF_buf1), .C(_2930__bF_buf7), .D(_2743_), .Y(_1316_) );
	INVX1 INVX1_1023 ( .A(micro_hash_synth_1_W_13__7_), .Y(_2745_) );
	INVX1 INVX1_1024 ( .A(bloque_in_111_), .Y(_2746_) );
	OAI22X1 OAI22X1_423 ( .A(_2746_), .B(_2925__bF_buf0), .C(_2930__bF_buf6), .D(_2745_), .Y(_1318_) );
	OAI21X1 OAI21X1_1143 ( .A(_3039_), .B(micro_hash_synth_1_W_7__0_), .C(_2731_), .Y(_2747_) );
	AOI21X1 AOI21X1_802 ( .A(_3039_), .B(micro_hash_synth_1_W_7__0_), .C(_2747_), .Y(_2748_) );
	OAI22X1 OAI22X1_424 ( .A(_2925__bF_buf15), .B(_2748_), .C(_2930__bF_buf5), .D(_1673_), .Y(_1319_) );
	OAI21X1 OAI21X1_1144 ( .A(_3040_), .B(micro_hash_synth_1_W_7__1_), .C(_2733_), .Y(_2749_) );
	AOI21X1 AOI21X1_803 ( .A(_3040_), .B(micro_hash_synth_1_W_7__1_), .C(_2749_), .Y(_2750_) );
	OAI22X1 OAI22X1_425 ( .A(_2925__bF_buf14), .B(_2750_), .C(_2930__bF_buf4), .D(_1707_), .Y(_1320_) );
	OAI21X1 OAI21X1_1145 ( .A(_3041_), .B(micro_hash_synth_1_W_7__2_), .C(_2735_), .Y(_2751_) );
	AOI21X1 AOI21X1_804 ( .A(_3041_), .B(micro_hash_synth_1_W_7__2_), .C(_2751_), .Y(_2752_) );
	OAI22X1 OAI22X1_426 ( .A(_2925__bF_buf13), .B(_2752_), .C(_2930__bF_buf3), .D(_1808_), .Y(_1321_) );
	OAI21X1 OAI21X1_1146 ( .A(_3042_), .B(micro_hash_synth_1_W_7__3_), .C(_2737_), .Y(_2753_) );
	AOI21X1 AOI21X1_805 ( .A(_3042_), .B(micro_hash_synth_1_W_7__3_), .C(_2753_), .Y(_2754_) );
	OAI22X1 OAI22X1_427 ( .A(_2925__bF_buf12), .B(_2754_), .C(_2930__bF_buf2), .D(_1938_), .Y(_1322_) );
	OAI21X1 OAI21X1_1147 ( .A(_3043_), .B(micro_hash_synth_1_W_7__4_), .C(_2739_), .Y(_2755_) );
	AOI21X1 AOI21X1_806 ( .A(_3043_), .B(micro_hash_synth_1_W_7__4_), .C(_2755_), .Y(_2756_) );
	OAI22X1 OAI22X1_428 ( .A(_2925__bF_buf11), .B(_2756_), .C(_2930__bF_buf1), .D(_2035_), .Y(_1323_) );
	OAI21X1 OAI21X1_1148 ( .A(_3044_), .B(micro_hash_synth_1_W_7__5_), .C(_2741_), .Y(_2757_) );
	AOI21X1 AOI21X1_807 ( .A(_3044_), .B(micro_hash_synth_1_W_7__5_), .C(_2757_), .Y(_2758_) );
	OAI22X1 OAI22X1_429 ( .A(_2925__bF_buf10), .B(_2758_), .C(_2930__bF_buf0), .D(_2092_), .Y(_1324_) );
	OAI21X1 OAI21X1_1149 ( .A(_3045_), .B(micro_hash_synth_1_W_7__6_), .C(_2743_), .Y(_2759_) );
	AOI21X1 AOI21X1_808 ( .A(_3045_), .B(micro_hash_synth_1_W_7__6_), .C(_2759_), .Y(_2760_) );
	OAI22X1 OAI22X1_430 ( .A(_2925__bF_buf9), .B(_2760_), .C(_2930__bF_buf13), .D(_2175_), .Y(_1325_) );
	OAI21X1 OAI21X1_1150 ( .A(_3046_), .B(micro_hash_synth_1_W_7__7_), .C(_2745_), .Y(_2761_) );
	AOI21X1 AOI21X1_809 ( .A(_3046_), .B(micro_hash_synth_1_W_7__7_), .C(_2761_), .Y(_2762_) );
	OAI22X1 OAI22X1_431 ( .A(_2925__bF_buf8), .B(_2762_), .C(_2930__bF_buf12), .D(_2642_), .Y(_1326_) );
	INVX1 INVX1_1025 ( .A(bloque_in_8_), .Y(_2763_) );
	OAI22X1 OAI22X1_432 ( .A(_2763_), .B(_2925__bF_buf7), .C(_2930__bF_buf11), .D(_3023_), .Y(_1327_) );
	INVX1 INVX1_1026 ( .A(bloque_in_9_), .Y(_2764_) );
	OAI22X1 OAI22X1_433 ( .A(_2764_), .B(_2925__bF_buf6), .C(_2930__bF_buf10), .D(_3024_), .Y(_1328_) );
	INVX1 INVX1_1027 ( .A(bloque_in_10_), .Y(_2765_) );
	OAI22X1 OAI22X1_434 ( .A(_2765_), .B(_2925__bF_buf5), .C(_2930__bF_buf9), .D(_3025_), .Y(_1329_) );
	INVX1 INVX1_1028 ( .A(bloque_in_11_), .Y(_2766_) );
	OAI22X1 OAI22X1_435 ( .A(_2766_), .B(_2925__bF_buf4), .C(_2930__bF_buf8), .D(_3026_), .Y(_1330_) );
	INVX1 INVX1_1029 ( .A(bloque_in_12_), .Y(_2767_) );
	OAI22X1 OAI22X1_436 ( .A(_2767_), .B(_2925__bF_buf3), .C(_2930__bF_buf7), .D(_3027_), .Y(_1331_) );
	INVX1 INVX1_1030 ( .A(bloque_in_13_), .Y(_2768_) );
	OAI22X1 OAI22X1_437 ( .A(_2768_), .B(_2925__bF_buf2), .C(_2930__bF_buf6), .D(_3028_), .Y(_1332_) );
	INVX1 INVX1_1031 ( .A(bloque_in_14_), .Y(_2769_) );
	OAI22X1 OAI22X1_438 ( .A(_2769_), .B(_2925__bF_buf1), .C(_2930__bF_buf5), .D(_3029_), .Y(_1334_) );
	INVX1 INVX1_1032 ( .A(bloque_in_15_), .Y(_2770_) );
	OAI22X1 OAI22X1_439 ( .A(_2770_), .B(_2925__bF_buf0), .C(_2930__bF_buf4), .D(_3030_), .Y(_1335_) );
	INVX1 INVX1_1033 ( .A(bloque_in_80_), .Y(_2771_) );
	NAND2X1 NAND2X1_634 ( .A(micro_hash_synth_1_W_10__0_), .B(_2459__bF_buf5), .Y(_2772_) );
	OAI21X1 OAI21X1_1151 ( .A(_2771_), .B(_2925__bF_buf15), .C(_2772_), .Y(_1336_) );
	INVX1 INVX1_1034 ( .A(bloque_in_81_), .Y(_2773_) );
	OAI22X1 OAI22X1_440 ( .A(_2773_), .B(_2925__bF_buf14), .C(_2930__bF_buf3), .D(_1736_), .Y(_1337_) );
	INVX1 INVX1_1035 ( .A(bloque_in_82_), .Y(_2774_) );
	OAI22X1 OAI22X1_441 ( .A(_2774_), .B(_2925__bF_buf13), .C(_2930__bF_buf2), .D(_1836_), .Y(_1338_) );
	INVX1 INVX1_1036 ( .A(bloque_in_83_), .Y(_2775_) );
	OAI22X1 OAI22X1_442 ( .A(_2775_), .B(_2925__bF_buf12), .C(_2930__bF_buf1), .D(_1951_), .Y(_1339_) );
	INVX1 INVX1_1037 ( .A(bloque_in_84_), .Y(_2776_) );
	OAI22X1 OAI22X1_443 ( .A(_2776_), .B(_2925__bF_buf11), .C(_2930__bF_buf0), .D(_2017_), .Y(_1340_) );
	INVX1 INVX1_1038 ( .A(bloque_in_85_), .Y(_2777_) );
	OAI22X1 OAI22X1_444 ( .A(_2777_), .B(_2925__bF_buf10), .C(_2930__bF_buf13), .D(_2119_), .Y(_1341_) );
	INVX1 INVX1_1039 ( .A(bloque_in_86_), .Y(_2778_) );
	OAI22X1 OAI22X1_445 ( .A(_2778_), .B(_2925__bF_buf9), .C(_2930__bF_buf12), .D(_2205_), .Y(_1342_) );
	INVX1 INVX1_1040 ( .A(bloque_in_87_), .Y(_2779_) );
	OAI22X1 OAI22X1_446 ( .A(_2779_), .B(_2925__bF_buf8), .C(_2930__bF_buf11), .D(_2455_), .Y(_1343_) );
	INVX1 INVX1_1041 ( .A(bloque_in_88_), .Y(_2780_) );
	NAND2X1 NAND2X1_635 ( .A(micro_hash_synth_1_W_11__0_), .B(_2459__bF_buf4), .Y(_2781_) );
	OAI21X1 OAI21X1_1152 ( .A(_2780_), .B(_2925__bF_buf7), .C(_2781_), .Y(_1344_) );
	INVX1 INVX1_1042 ( .A(bloque_in_89_), .Y(_2782_) );
	OAI22X1 OAI22X1_447 ( .A(_2782_), .B(_2925__bF_buf6), .C(_2930__bF_buf10), .D(_2966_), .Y(_1345_) );
	INVX1 INVX1_1043 ( .A(bloque_in_90_), .Y(_2783_) );
	OAI22X1 OAI22X1_448 ( .A(_2783_), .B(_2925__bF_buf5), .C(_2930__bF_buf9), .D(_2971_), .Y(_1346_) );
	INVX1 INVX1_1044 ( .A(bloque_in_91_), .Y(_2784_) );
	NAND2X1 NAND2X1_636 ( .A(micro_hash_synth_1_W_11__3_), .B(_2459__bF_buf3), .Y(_2785_) );
	OAI21X1 OAI21X1_1153 ( .A(_2784_), .B(_2925__bF_buf4), .C(_2785_), .Y(_1347_) );
	INVX1 INVX1_1045 ( .A(bloque_in_92_), .Y(_2786_) );
	NAND2X1 NAND2X1_637 ( .A(micro_hash_synth_1_W_11__4_), .B(_2459__bF_buf2), .Y(_2787_) );
	OAI21X1 OAI21X1_1154 ( .A(_2786_), .B(_2925__bF_buf3), .C(_2787_), .Y(_1348_) );
	INVX1 INVX1_1046 ( .A(bloque_in_93_), .Y(_2788_) );
	NAND2X1 NAND2X1_638 ( .A(micro_hash_synth_1_W_11__5_), .B(_2459__bF_buf1), .Y(_2789_) );
	OAI21X1 OAI21X1_1155 ( .A(_2788_), .B(_2925__bF_buf2), .C(_2789_), .Y(_1349_) );
	INVX1 INVX1_1047 ( .A(bloque_in_94_), .Y(_2790_) );
	NAND2X1 NAND2X1_639 ( .A(micro_hash_synth_1_W_11__6_), .B(_2459__bF_buf0), .Y(_2791_) );
	OAI21X1 OAI21X1_1156 ( .A(_2790_), .B(_2925__bF_buf1), .C(_2791_), .Y(_1350_) );
	INVX1 INVX1_1048 ( .A(bloque_in_95_), .Y(_2792_) );
	NAND2X1 NAND2X1_640 ( .A(micro_hash_synth_1_W_11__7_), .B(_2459__bF_buf6), .Y(_2793_) );
	OAI21X1 OAI21X1_1157 ( .A(_2792_), .B(_2925__bF_buf0), .C(_2793_), .Y(_1351_) );
	INVX1 INVX1_1049 ( .A(bloque_in_16_), .Y(_2794_) );
	OAI22X1 OAI22X1_449 ( .A(_2794_), .B(_2925__bF_buf15), .C(_2930__bF_buf8), .D(_3039_), .Y(_1352_) );
	INVX1 INVX1_1050 ( .A(bloque_in_17_), .Y(_2795_) );
	OAI22X1 OAI22X1_450 ( .A(_2795_), .B(_2925__bF_buf14), .C(_2930__bF_buf7), .D(_3040_), .Y(_1353_) );
	INVX1 INVX1_1051 ( .A(bloque_in_18_), .Y(_2796_) );
	OAI22X1 OAI22X1_451 ( .A(_2796_), .B(_2925__bF_buf13), .C(_2930__bF_buf6), .D(_3041_), .Y(_1354_) );
	INVX1 INVX1_1052 ( .A(bloque_in_19_), .Y(_2797_) );
	OAI22X1 OAI22X1_452 ( .A(_2797_), .B(_2925__bF_buf12), .C(_2930__bF_buf5), .D(_3042_), .Y(_1355_) );
	INVX1 INVX1_1053 ( .A(bloque_in_20_), .Y(_2798_) );
	OAI22X1 OAI22X1_453 ( .A(_2798_), .B(_2925__bF_buf11), .C(_2930__bF_buf4), .D(_3043_), .Y(_1356_) );
	INVX1 INVX1_1054 ( .A(bloque_in_21_), .Y(_2799_) );
	OAI22X1 OAI22X1_454 ( .A(_2799_), .B(_2925__bF_buf10), .C(_2930__bF_buf3), .D(_3044_), .Y(_1357_) );
	INVX1 INVX1_1055 ( .A(bloque_in_22_), .Y(_2800_) );
	OAI22X1 OAI22X1_455 ( .A(_2800_), .B(_2925__bF_buf9), .C(_2930__bF_buf2), .D(_3045_), .Y(_1358_) );
	INVX1 INVX1_1056 ( .A(bloque_in_23_), .Y(_2801_) );
	OAI22X1 OAI22X1_456 ( .A(_2801_), .B(_2925__bF_buf8), .C(_2930__bF_buf1), .D(_3046_), .Y(_1359_) );
	INVX1 INVX1_1057 ( .A(micro_hash_synth_1_W_27__0_), .Y(_2802_) );
	OAI21X1 OAI21X1_1158 ( .A(_2731_), .B(micro_hash_synth_1_W_18__0_), .C(_2434_), .Y(_2803_) );
	AOI21X1 AOI21X1_810 ( .A(_2731_), .B(micro_hash_synth_1_W_18__0_), .C(_2803_), .Y(_2804_) );
	OAI22X1 OAI22X1_457 ( .A(_2925__bF_buf7), .B(_2804_), .C(_2930__bF_buf0), .D(_2802_), .Y(_1360_) );
	INVX1 INVX1_1058 ( .A(micro_hash_synth_1_W_27__1_), .Y(_2805_) );
	OAI21X1 OAI21X1_1159 ( .A(_2733_), .B(micro_hash_synth_1_W_18__1_), .C(_1723_), .Y(_2806_) );
	AOI21X1 AOI21X1_811 ( .A(_2733_), .B(micro_hash_synth_1_W_18__1_), .C(_2806_), .Y(_2807_) );
	OAI22X1 OAI22X1_458 ( .A(_2925__bF_buf6), .B(_2807_), .C(_2930__bF_buf13), .D(_2805_), .Y(_1361_) );
	INVX1 INVX1_1059 ( .A(micro_hash_synth_1_W_27__2_), .Y(_2808_) );
	OAI21X1 OAI21X1_1160 ( .A(_2735_), .B(micro_hash_synth_1_W_18__2_), .C(_1819_), .Y(_2809_) );
	AOI21X1 AOI21X1_812 ( .A(_2735_), .B(micro_hash_synth_1_W_18__2_), .C(_2809_), .Y(_2810_) );
	OAI22X1 OAI22X1_459 ( .A(_2925__bF_buf5), .B(_2810_), .C(_2930__bF_buf12), .D(_2808_), .Y(_1362_) );
	INVX1 INVX1_1060 ( .A(micro_hash_synth_1_W_27__3_), .Y(_2811_) );
	OAI21X1 OAI21X1_1161 ( .A(_2737_), .B(micro_hash_synth_1_W_18__3_), .C(_1919_), .Y(_2812_) );
	AOI21X1 AOI21X1_813 ( .A(_2737_), .B(micro_hash_synth_1_W_18__3_), .C(_2812_), .Y(_2813_) );
	OAI22X1 OAI22X1_460 ( .A(_2925__bF_buf4), .B(_2813_), .C(_2930__bF_buf11), .D(_2811_), .Y(_1363_) );
	INVX1 INVX1_1061 ( .A(micro_hash_synth_1_W_27__4_), .Y(_2814_) );
	OAI21X1 OAI21X1_1162 ( .A(_2739_), .B(micro_hash_synth_1_W_18__4_), .C(_2003_), .Y(_2815_) );
	AOI21X1 AOI21X1_814 ( .A(_2739_), .B(micro_hash_synth_1_W_18__4_), .C(_2815_), .Y(_2816_) );
	OAI22X1 OAI22X1_461 ( .A(_2925__bF_buf3), .B(_2816_), .C(_2930__bF_buf10), .D(_2814_), .Y(_1364_) );
	INVX1 INVX1_1062 ( .A(micro_hash_synth_1_W_27__5_), .Y(_2817_) );
	OAI21X1 OAI21X1_1163 ( .A(_2741_), .B(micro_hash_synth_1_W_18__5_), .C(_2105_), .Y(_2818_) );
	AOI21X1 AOI21X1_815 ( .A(_2741_), .B(micro_hash_synth_1_W_18__5_), .C(_2818_), .Y(_2819_) );
	OAI22X1 OAI22X1_462 ( .A(_2925__bF_buf2), .B(_2819_), .C(_2930__bF_buf9), .D(_2817_), .Y(_1365_) );
	INVX1 INVX1_1063 ( .A(micro_hash_synth_1_W_27__6_), .Y(_2820_) );
	OAI21X1 OAI21X1_1164 ( .A(_2743_), .B(micro_hash_synth_1_W_18__6_), .C(_2186_), .Y(_2821_) );
	AOI21X1 AOI21X1_816 ( .A(_2743_), .B(micro_hash_synth_1_W_18__6_), .C(_2821_), .Y(_2822_) );
	OAI22X1 OAI22X1_463 ( .A(_2925__bF_buf1), .B(_2822_), .C(_2930__bF_buf8), .D(_2820_), .Y(_1366_) );
	INVX1 INVX1_1064 ( .A(micro_hash_synth_1_W_27__7_), .Y(_2823_) );
	OAI21X1 OAI21X1_1165 ( .A(_2745_), .B(micro_hash_synth_1_W_18__7_), .C(_2258_), .Y(_2824_) );
	AOI21X1 AOI21X1_817 ( .A(_2745_), .B(micro_hash_synth_1_W_18__7_), .C(_2824_), .Y(_2825_) );
	OAI22X1 OAI22X1_464 ( .A(_2925__bF_buf0), .B(_2825_), .C(_2930__bF_buf7), .D(_2823_), .Y(_1367_) );
	INVX1 INVX1_1065 ( .A(micro_hash_synth_1_W_28__0_), .Y(_2826_) );
	OAI21X1 OAI21X1_1166 ( .A(_2653_), .B(micro_hash_synth_1_W_19__0_), .C(_2962_), .Y(_2827_) );
	AOI21X1 AOI21X1_818 ( .A(_2653_), .B(micro_hash_synth_1_W_19__0_), .C(_2827_), .Y(_2828_) );
	OAI22X1 OAI22X1_465 ( .A(_2925__bF_buf15), .B(_2828_), .C(_2930__bF_buf6), .D(_2826_), .Y(_1368_) );
	INVX1 INVX1_1066 ( .A(micro_hash_synth_1_W_28__1_), .Y(_2829_) );
	OAI21X1 OAI21X1_1167 ( .A(_2655_), .B(micro_hash_synth_1_W_19__1_), .C(_2965_), .Y(_2830_) );
	AOI21X1 AOI21X1_819 ( .A(_2655_), .B(micro_hash_synth_1_W_19__1_), .C(_2830_), .Y(_2831_) );
	OAI22X1 OAI22X1_466 ( .A(_2925__bF_buf14), .B(_2831_), .C(_2930__bF_buf5), .D(_2829_), .Y(_1369_) );
	INVX1 INVX1_1067 ( .A(micro_hash_synth_1_W_28__2_), .Y(_2832_) );
	OAI21X1 OAI21X1_1168 ( .A(_2657_), .B(micro_hash_synth_1_W_19__2_), .C(_2970_), .Y(_2833_) );
	AOI21X1 AOI21X1_820 ( .A(_2657_), .B(micro_hash_synth_1_W_19__2_), .C(_2833_), .Y(_2834_) );
	OAI22X1 OAI22X1_467 ( .A(_2925__bF_buf13), .B(_2834_), .C(_2930__bF_buf4), .D(_2832_), .Y(_1370_) );
	INVX1 INVX1_1068 ( .A(micro_hash_synth_1_W_28__3_), .Y(_2835_) );
	OAI21X1 OAI21X1_1169 ( .A(_2659_), .B(micro_hash_synth_1_W_19__3_), .C(_2975_), .Y(_2836_) );
	AOI21X1 AOI21X1_821 ( .A(_2659_), .B(micro_hash_synth_1_W_19__3_), .C(_2836_), .Y(_2837_) );
	OAI22X1 OAI22X1_468 ( .A(_2925__bF_buf12), .B(_2837_), .C(_2930__bF_buf3), .D(_2835_), .Y(_1371_) );
	INVX1 INVX1_1069 ( .A(micro_hash_synth_1_W_28__4_), .Y(_2838_) );
	OAI21X1 OAI21X1_1170 ( .A(_2661_), .B(micro_hash_synth_1_W_19__4_), .C(_2978_), .Y(_2839_) );
	AOI21X1 AOI21X1_822 ( .A(_2661_), .B(micro_hash_synth_1_W_19__4_), .C(_2839_), .Y(_2840_) );
	OAI22X1 OAI22X1_469 ( .A(_2925__bF_buf11), .B(_2840_), .C(_2930__bF_buf2), .D(_2838_), .Y(_1372_) );
	INVX1 INVX1_1070 ( .A(micro_hash_synth_1_W_28__5_), .Y(_2841_) );
	OAI21X1 OAI21X1_1171 ( .A(_2663_), .B(micro_hash_synth_1_W_19__5_), .C(_2981_), .Y(_2842_) );
	AOI21X1 AOI21X1_823 ( .A(_2663_), .B(micro_hash_synth_1_W_19__5_), .C(_2842_), .Y(_2843_) );
	OAI22X1 OAI22X1_470 ( .A(_2925__bF_buf10), .B(_2843_), .C(_2930__bF_buf1), .D(_2841_), .Y(_1373_) );
	INVX1 INVX1_1071 ( .A(micro_hash_synth_1_W_28__6_), .Y(_2844_) );
	OAI21X1 OAI21X1_1172 ( .A(_2665_), .B(micro_hash_synth_1_W_19__6_), .C(_2984_), .Y(_2845_) );
	AOI21X1 AOI21X1_824 ( .A(_2665_), .B(micro_hash_synth_1_W_19__6_), .C(_2845_), .Y(_2846_) );
	OAI22X1 OAI22X1_471 ( .A(_2925__bF_buf9), .B(_2846_), .C(_2930__bF_buf0), .D(_2844_), .Y(_1374_) );
	INVX1 INVX1_1072 ( .A(micro_hash_synth_1_W_28__7_), .Y(_2847_) );
	OAI21X1 OAI21X1_1173 ( .A(_2667_), .B(micro_hash_synth_1_W_19__7_), .C(_2987_), .Y(_2848_) );
	AOI21X1 AOI21X1_825 ( .A(_2667_), .B(micro_hash_synth_1_W_19__7_), .C(_2848_), .Y(_2849_) );
	OAI22X1 OAI22X1_472 ( .A(_2925__bF_buf8), .B(_2849_), .C(_2930__bF_buf13), .D(_2847_), .Y(_1375_) );
	NAND2X1 NAND2X1_641 ( .A(micro_hash_synth_1_W_29__0_), .B(_2459__bF_buf5), .Y(_2850_) );
	OAI21X1 OAI21X1_1174 ( .A(_2677_), .B(micro_hash_synth_1_W_20__0_), .C(_2918_), .Y(_2851_) );
	AOI21X1 AOI21X1_826 ( .A(_2677_), .B(micro_hash_synth_1_W_20__0_), .C(_2851_), .Y(_2852_) );
	OAI21X1 OAI21X1_1175 ( .A(_2925__bF_buf7), .B(_2852_), .C(_2850_), .Y(_1376_) );
	OAI21X1 OAI21X1_1176 ( .A(_2680_), .B(micro_hash_synth_1_W_20__1_), .C(_2933_), .Y(_2853_) );
	AOI21X1 AOI21X1_827 ( .A(_2680_), .B(micro_hash_synth_1_W_20__1_), .C(_2853_), .Y(_2854_) );
	OAI22X1 OAI22X1_473 ( .A(_2925__bF_buf6), .B(_2854_), .C(_2930__bF_buf12), .D(_1714_), .Y(_1377_) );
	OAI21X1 OAI21X1_1177 ( .A(_2683_), .B(micro_hash_synth_1_W_20__2_), .C(_2938_), .Y(_2855_) );
	AOI21X1 AOI21X1_828 ( .A(_2683_), .B(micro_hash_synth_1_W_20__2_), .C(_2855_), .Y(_2856_) );
	OAI22X1 OAI22X1_474 ( .A(_2925__bF_buf5), .B(_2856_), .C(_2930__bF_buf11), .D(_1864_), .Y(_1378_) );
	NAND2X1 NAND2X1_642 ( .A(micro_hash_synth_1_W_29__3_), .B(_2459__bF_buf4), .Y(_2857_) );
	OAI21X1 OAI21X1_1178 ( .A(_2686_), .B(micro_hash_synth_1_W_20__3_), .C(_2943_), .Y(_2858_) );
	AOI21X1 AOI21X1_829 ( .A(_2686_), .B(micro_hash_synth_1_W_20__3_), .C(_2858_), .Y(_2859_) );
	OAI21X1 OAI21X1_1179 ( .A(_2925__bF_buf4), .B(_2859_), .C(_2857_), .Y(_1379_) );
	NAND2X1 NAND2X1_643 ( .A(micro_hash_synth_1_W_29__4_), .B(_2459__bF_buf3), .Y(_2860_) );
	OAI21X1 OAI21X1_1180 ( .A(_2689_), .B(micro_hash_synth_1_W_20__4_), .C(_2946_), .Y(_2861_) );
	AOI21X1 AOI21X1_830 ( .A(_2689_), .B(micro_hash_synth_1_W_20__4_), .C(_2861_), .Y(_2862_) );
	OAI21X1 OAI21X1_1181 ( .A(_2925__bF_buf3), .B(_2862_), .C(_2860_), .Y(_1380_) );
	NAND2X1 NAND2X1_644 ( .A(micro_hash_synth_1_W_29__5_), .B(_2459__bF_buf2), .Y(_2863_) );
	OAI21X1 OAI21X1_1182 ( .A(_2692_), .B(micro_hash_synth_1_W_20__5_), .C(_2949_), .Y(_2864_) );
	AOI21X1 AOI21X1_831 ( .A(_2692_), .B(micro_hash_synth_1_W_20__5_), .C(_2864_), .Y(_2865_) );
	OAI21X1 OAI21X1_1183 ( .A(_2925__bF_buf2), .B(_2865_), .C(_2863_), .Y(_1381_) );
	NAND2X1 NAND2X1_645 ( .A(micro_hash_synth_1_W_29__6_), .B(_2459__bF_buf1), .Y(_2866_) );
	OAI21X1 OAI21X1_1184 ( .A(_2197_), .B(micro_hash_synth_1_W_20__6_), .C(_2952_), .Y(_2867_) );
	AOI21X1 AOI21X1_832 ( .A(_2197_), .B(micro_hash_synth_1_W_20__6_), .C(_2867_), .Y(_2868_) );
	OAI21X1 OAI21X1_1185 ( .A(_2925__bF_buf1), .B(_2868_), .C(_2866_), .Y(_1382_) );
	NAND2X1 NAND2X1_646 ( .A(micro_hash_synth_1_W_29__7_), .B(_2459__bF_buf0), .Y(_2869_) );
	OAI21X1 OAI21X1_1186 ( .A(_2266_), .B(micro_hash_synth_1_W_20__7_), .C(_2957_), .Y(_2870_) );
	AOI21X1 AOI21X1_833 ( .A(_2266_), .B(micro_hash_synth_1_W_20__7_), .C(_2870_), .Y(_2871_) );
	OAI21X1 OAI21X1_1187 ( .A(_2925__bF_buf0), .B(_2871_), .C(_2869_), .Y(_1383_) );
	NAND2X1 NAND2X1_647 ( .A(micro_hash_synth_1_W_30__0_), .B(_2459__bF_buf6), .Y(_2872_) );
	OAI21X1 OAI21X1_1188 ( .A(_1673_), .B(micro_hash_synth_1_W_21__0_), .C(_2802_), .Y(_2873_) );
	AOI21X1 AOI21X1_834 ( .A(_1673_), .B(micro_hash_synth_1_W_21__0_), .C(_2873_), .Y(_2874_) );
	OAI21X1 OAI21X1_1189 ( .A(_2925__bF_buf15), .B(_2874_), .C(_2872_), .Y(_1384_) );
	NAND2X1 NAND2X1_648 ( .A(micro_hash_synth_1_W_30__1_), .B(_2459__bF_buf5), .Y(_2875_) );
	OAI21X1 OAI21X1_1190 ( .A(_1707_), .B(micro_hash_synth_1_W_21__1_), .C(_2805_), .Y(_2876_) );
	AOI21X1 AOI21X1_835 ( .A(_1707_), .B(micro_hash_synth_1_W_21__1_), .C(_2876_), .Y(_2877_) );
	OAI21X1 OAI21X1_1191 ( .A(_2925__bF_buf14), .B(_2877_), .C(_2875_), .Y(_1385_) );
	NAND2X1 NAND2X1_649 ( .A(micro_hash_synth_1_W_30__2_), .B(_2459__bF_buf4), .Y(_2878_) );
	OAI21X1 OAI21X1_1192 ( .A(_1808_), .B(micro_hash_synth_1_W_21__2_), .C(_2808_), .Y(_2879_) );
	AOI21X1 AOI21X1_836 ( .A(_1808_), .B(micro_hash_synth_1_W_21__2_), .C(_2879_), .Y(_2880_) );
	OAI21X1 OAI21X1_1193 ( .A(_2925__bF_buf13), .B(_2880_), .C(_2878_), .Y(_1386_) );
	NAND2X1 NAND2X1_650 ( .A(micro_hash_synth_1_W_30__3_), .B(_2459__bF_buf3), .Y(_2881_) );
	OAI21X1 OAI21X1_1194 ( .A(_1938_), .B(micro_hash_synth_1_W_21__3_), .C(_2811_), .Y(_2882_) );
	AOI21X1 AOI21X1_837 ( .A(_1938_), .B(micro_hash_synth_1_W_21__3_), .C(_2882_), .Y(_2883_) );
	OAI21X1 OAI21X1_1195 ( .A(_2925__bF_buf12), .B(_2883_), .C(_2881_), .Y(_1387_) );
	NAND2X1 NAND2X1_651 ( .A(micro_hash_synth_1_W_30__4_), .B(_2459__bF_buf2), .Y(_2884_) );
	OAI21X1 OAI21X1_1196 ( .A(_2035_), .B(micro_hash_synth_1_W_21__4_), .C(_2814_), .Y(_2885_) );
	AOI21X1 AOI21X1_838 ( .A(_2035_), .B(micro_hash_synth_1_W_21__4_), .C(_2885_), .Y(_2886_) );
	OAI21X1 OAI21X1_1197 ( .A(_2925__bF_buf11), .B(_2886_), .C(_2884_), .Y(_1388_) );
	NAND2X1 NAND2X1_652 ( .A(micro_hash_synth_1_W_30__5_), .B(_2459__bF_buf1), .Y(_2887_) );
	OAI21X1 OAI21X1_1198 ( .A(_2092_), .B(micro_hash_synth_1_W_21__5_), .C(_2817_), .Y(_2888_) );
	AOI21X1 AOI21X1_839 ( .A(_2092_), .B(micro_hash_synth_1_W_21__5_), .C(_2888_), .Y(_2889_) );
	OAI21X1 OAI21X1_1199 ( .A(_2925__bF_buf10), .B(_2889_), .C(_2887_), .Y(_1389_) );
	NAND2X1 NAND2X1_653 ( .A(micro_hash_synth_1_W_30__6_), .B(_2459__bF_buf0), .Y(_2890_) );
	OAI21X1 OAI21X1_1200 ( .A(_2175_), .B(micro_hash_synth_1_W_21__6_), .C(_2820_), .Y(_2891_) );
	AOI21X1 AOI21X1_840 ( .A(_2175_), .B(micro_hash_synth_1_W_21__6_), .C(_2891_), .Y(_2892_) );
	OAI21X1 OAI21X1_1201 ( .A(_2925__bF_buf9), .B(_2892_), .C(_2890_), .Y(_1390_) );
	NAND2X1 NAND2X1_654 ( .A(micro_hash_synth_1_W_30__7_), .B(_2459__bF_buf6), .Y(_2893_) );
	OAI21X1 OAI21X1_1202 ( .A(_2642_), .B(micro_hash_synth_1_W_21__7_), .C(_2823_), .Y(_2894_) );
	AOI21X1 AOI21X1_841 ( .A(_2642_), .B(micro_hash_synth_1_W_21__7_), .C(_2894_), .Y(_2895_) );
	OAI21X1 OAI21X1_1203 ( .A(_2925__bF_buf8), .B(_2895_), .C(_2893_), .Y(_1391_) );
	NAND2X1 NAND2X1_655 ( .A(micro_hash_synth_1_W_31__0_), .B(_2459__bF_buf5), .Y(_2896_) );
	OAI21X1 OAI21X1_1204 ( .A(_2574_), .B(micro_hash_synth_1_W_22__0_), .C(_2826_), .Y(_2897_) );
	AOI21X1 AOI21X1_842 ( .A(_2574_), .B(micro_hash_synth_1_W_22__0_), .C(_2897_), .Y(_2898_) );
	OAI21X1 OAI21X1_1205 ( .A(_2925__bF_buf7), .B(_2898_), .C(_2896_), .Y(_1392_) );
	OAI21X1 OAI21X1_1206 ( .A(_2579_), .B(micro_hash_synth_1_W_22__1_), .C(_2829_), .Y(_2899_) );
	AOI21X1 AOI21X1_843 ( .A(_2579_), .B(micro_hash_synth_1_W_22__1_), .C(_2899_), .Y(_2900_) );
	OAI22X1 OAI22X1_475 ( .A(_2925__bF_buf6), .B(_2900_), .C(_2930__bF_buf10), .D(_1719_), .Y(_1393_) );
	OAI21X1 OAI21X1_1207 ( .A(_2584_), .B(micro_hash_synth_1_W_22__2_), .C(_2832_), .Y(_2901_) );
	AOI21X1 AOI21X1_844 ( .A(_2584_), .B(micro_hash_synth_1_W_22__2_), .C(_2901_), .Y(_2902_) );
	OAI22X1 OAI22X1_476 ( .A(_2925__bF_buf5), .B(_2902_), .C(_2930__bF_buf9), .D(_1869_), .Y(_1394_) );
	NAND2X1 NAND2X1_656 ( .A(micro_hash_synth_1_W_31__3_), .B(_2459__bF_buf4), .Y(_2903_) );
	OAI21X1 OAI21X1_1208 ( .A(_2589_), .B(micro_hash_synth_1_W_22__3_), .C(_2835_), .Y(_2904_) );
	AOI21X1 AOI21X1_845 ( .A(_2589_), .B(micro_hash_synth_1_W_22__3_), .C(_2904_), .Y(_2905_) );
	OAI21X1 OAI21X1_1209 ( .A(_2925__bF_buf4), .B(_2905_), .C(_2903_), .Y(_1395_) );
	NAND2X1 NAND2X1_657 ( .A(micro_hash_synth_1_W_31__4_), .B(_2459__bF_buf3), .Y(_2906_) );
	OAI21X1 OAI21X1_1210 ( .A(_2594_), .B(micro_hash_synth_1_W_22__4_), .C(_2838_), .Y(_2907_) );
	AOI21X1 AOI21X1_846 ( .A(_2594_), .B(micro_hash_synth_1_W_22__4_), .C(_2907_), .Y(_2908_) );
	OAI21X1 OAI21X1_1211 ( .A(_2925__bF_buf3), .B(_2908_), .C(_2906_), .Y(_1396_) );
	NAND2X1 NAND2X1_658 ( .A(micro_hash_synth_1_W_31__5_), .B(_2459__bF_buf2), .Y(_2909_) );
	OAI21X1 OAI21X1_1212 ( .A(_2599_), .B(micro_hash_synth_1_W_22__5_), .C(_2841_), .Y(_2910_) );
	AOI21X1 AOI21X1_847 ( .A(_2599_), .B(micro_hash_synth_1_W_22__5_), .C(_2910_), .Y(_2911_) );
	OAI21X1 OAI21X1_1213 ( .A(_2925__bF_buf2), .B(_2911_), .C(_2909_), .Y(_1397_) );
	NAND2X1 NAND2X1_659 ( .A(micro_hash_synth_1_W_31__6_), .B(_2459__bF_buf1), .Y(_2912_) );
	OAI21X1 OAI21X1_1214 ( .A(_2603_), .B(micro_hash_synth_1_W_22__6_), .C(_2844_), .Y(_2913_) );
	AOI21X1 AOI21X1_848 ( .A(_2603_), .B(micro_hash_synth_1_W_22__6_), .C(_2913_), .Y(_2914_) );
	OAI21X1 OAI21X1_1215 ( .A(_2925__bF_buf1), .B(_2914_), .C(_2912_), .Y(_1398_) );
	NAND2X1 NAND2X1_660 ( .A(micro_hash_synth_1_W_31__7_), .B(_2459__bF_buf0), .Y(_2915_) );
	OAI21X1 OAI21X1_1216 ( .A(_2607_), .B(micro_hash_synth_1_W_22__7_), .C(_2847_), .Y(_2916_) );
	AOI21X1 AOI21X1_849 ( .A(_2607_), .B(micro_hash_synth_1_W_22__7_), .C(_2916_), .Y(_2917_) );
	OAI21X1 OAI21X1_1217 ( .A(_2925__bF_buf0), .B(_2917_), .C(_2915_), .Y(_1399_) );
	DFFPOSX1 DFFPOSX1_879 ( .CLK(clk_bF_buf33), .D(_1432_), .Q(micro_hash_synth_1_W_22__0_) );
	DFFPOSX1 DFFPOSX1_880 ( .CLK(clk_bF_buf32), .D(_1433_), .Q(micro_hash_synth_1_W_22__1_) );
	DFFPOSX1 DFFPOSX1_881 ( .CLK(clk_bF_buf31), .D(_1435_), .Q(micro_hash_synth_1_W_22__2_) );
	DFFPOSX1 DFFPOSX1_882 ( .CLK(clk_bF_buf30), .D(_1436_), .Q(micro_hash_synth_1_W_22__3_) );
	DFFPOSX1 DFFPOSX1_883 ( .CLK(clk_bF_buf29), .D(_1437_), .Q(micro_hash_synth_1_W_22__4_) );
	DFFPOSX1 DFFPOSX1_884 ( .CLK(clk_bF_buf28), .D(_1438_), .Q(micro_hash_synth_1_W_22__5_) );
	DFFPOSX1 DFFPOSX1_885 ( .CLK(clk_bF_buf27), .D(_1439_), .Q(micro_hash_synth_1_W_22__6_) );
	DFFPOSX1 DFFPOSX1_886 ( .CLK(clk_bF_buf26), .D(_1440_), .Q(micro_hash_synth_1_W_22__7_) );
	DFFPOSX1 DFFPOSX1_887 ( .CLK(clk_bF_buf25), .D(_1267_), .Q(micro_hash_synth_1_W_0__0_) );
	DFFPOSX1 DFFPOSX1_888 ( .CLK(clk_bF_buf24), .D(_1268_), .Q(micro_hash_synth_1_W_0__1_) );
	DFFPOSX1 DFFPOSX1_889 ( .CLK(clk_bF_buf23), .D(_1270_), .Q(micro_hash_synth_1_W_0__2_) );
	DFFPOSX1 DFFPOSX1_890 ( .CLK(clk_bF_buf22), .D(_1271_), .Q(micro_hash_synth_1_W_0__3_) );
	DFFPOSX1 DFFPOSX1_891 ( .CLK(clk_bF_buf21), .D(_1272_), .Q(micro_hash_synth_1_W_0__4_) );
	DFFPOSX1 DFFPOSX1_892 ( .CLK(clk_bF_buf20), .D(_1273_), .Q(micro_hash_synth_1_W_0__5_) );
	DFFPOSX1 DFFPOSX1_893 ( .CLK(clk_bF_buf19), .D(_1274_), .Q(micro_hash_synth_1_W_0__6_) );
	DFFPOSX1 DFFPOSX1_894 ( .CLK(clk_bF_buf18), .D(_1275_), .Q(micro_hash_synth_1_W_0__7_) );
	DFFPOSX1 DFFPOSX1_895 ( .CLK(clk_bF_buf17), .D(_1488_), .Q(micro_hash_synth_1_W_19__0_) );
	DFFPOSX1 DFFPOSX1_896 ( .CLK(clk_bF_buf16), .D(_1489_), .Q(micro_hash_synth_1_W_19__1_) );
	DFFPOSX1 DFFPOSX1_897 ( .CLK(clk_bF_buf15), .D(_1490_), .Q(micro_hash_synth_1_W_19__2_) );
	DFFPOSX1 DFFPOSX1_898 ( .CLK(clk_bF_buf14), .D(_1491_), .Q(micro_hash_synth_1_W_19__3_) );
	DFFPOSX1 DFFPOSX1_899 ( .CLK(clk_bF_buf13), .D(_1493_), .Q(micro_hash_synth_1_W_19__4_) );
	DFFPOSX1 DFFPOSX1_900 ( .CLK(clk_bF_buf12), .D(_1494_), .Q(micro_hash_synth_1_W_19__5_) );
	DFFPOSX1 DFFPOSX1_901 ( .CLK(clk_bF_buf11), .D(_1495_), .Q(micro_hash_synth_1_W_19__6_) );
	DFFPOSX1 DFFPOSX1_902 ( .CLK(clk_bF_buf10), .D(_1496_), .Q(micro_hash_synth_1_W_19__7_) );
	DFFPOSX1 DFFPOSX1_903 ( .CLK(clk_bF_buf9), .D(_1468_), .Q(micro_hash_synth_1_W_20__0_) );
	DFFPOSX1 DFFPOSX1_904 ( .CLK(clk_bF_buf8), .D(_1469_), .Q(micro_hash_synth_1_W_20__1_) );
	DFFPOSX1 DFFPOSX1_905 ( .CLK(clk_bF_buf7), .D(_1470_), .Q(micro_hash_synth_1_W_20__2_) );
	DFFPOSX1 DFFPOSX1_906 ( .CLK(clk_bF_buf6), .D(_1471_), .Q(micro_hash_synth_1_W_20__3_) );
	DFFPOSX1 DFFPOSX1_907 ( .CLK(clk_bF_buf5), .D(_1472_), .Q(micro_hash_synth_1_W_20__4_) );
	DFFPOSX1 DFFPOSX1_908 ( .CLK(clk_bF_buf4), .D(_1473_), .Q(micro_hash_synth_1_W_20__5_) );
	DFFPOSX1 DFFPOSX1_909 ( .CLK(clk_bF_buf3), .D(_1474_), .Q(micro_hash_synth_1_W_20__6_) );
	DFFPOSX1 DFFPOSX1_910 ( .CLK(clk_bF_buf2), .D(_1475_), .Q(micro_hash_synth_1_W_20__7_) );
	DFFPOSX1 DFFPOSX1_911 ( .CLK(clk_bF_buf1), .D(_1459_), .Q(micro_hash_synth_1_W_21__0_) );
	DFFPOSX1 DFFPOSX1_912 ( .CLK(clk_bF_buf0), .D(_1460_), .Q(micro_hash_synth_1_W_21__1_) );
	DFFPOSX1 DFFPOSX1_913 ( .CLK(clk_bF_buf113), .D(_1461_), .Q(micro_hash_synth_1_W_21__2_) );
	DFFPOSX1 DFFPOSX1_914 ( .CLK(clk_bF_buf112), .D(_1462_), .Q(micro_hash_synth_1_W_21__3_) );
	DFFPOSX1 DFFPOSX1_915 ( .CLK(clk_bF_buf111), .D(_1463_), .Q(micro_hash_synth_1_W_21__4_) );
	DFFPOSX1 DFFPOSX1_916 ( .CLK(clk_bF_buf110), .D(_1464_), .Q(micro_hash_synth_1_W_21__5_) );
	DFFPOSX1 DFFPOSX1_917 ( .CLK(clk_bF_buf109), .D(_1465_), .Q(micro_hash_synth_1_W_21__6_) );
	DFFPOSX1 DFFPOSX1_918 ( .CLK(clk_bF_buf108), .D(_1466_), .Q(micro_hash_synth_1_W_21__7_) );
	DFFPOSX1 DFFPOSX1_919 ( .CLK(clk_bF_buf107), .D(_1237__0_), .Q(Hhash_synth1_0_) );
	DFFPOSX1 DFFPOSX1_920 ( .CLK(clk_bF_buf106), .D(_1237__1_), .Q(Hhash_synth1_1_) );
	DFFPOSX1 DFFPOSX1_921 ( .CLK(clk_bF_buf105), .D(_1237__2_), .Q(Hhash_synth1_2_) );
	DFFPOSX1 DFFPOSX1_922 ( .CLK(clk_bF_buf104), .D(_1237__3_), .Q(Hhash_synth1_3_) );
	DFFPOSX1 DFFPOSX1_923 ( .CLK(clk_bF_buf103), .D(_1237__4_), .Q(Hhash_synth1_4_) );
	DFFPOSX1 DFFPOSX1_924 ( .CLK(clk_bF_buf102), .D(_1237__5_), .Q(Hhash_synth1_5_) );
	DFFPOSX1 DFFPOSX1_925 ( .CLK(clk_bF_buf101), .D(_1237__6_), .Q(Hhash_synth1_6_) );
	DFFPOSX1 DFFPOSX1_926 ( .CLK(clk_bF_buf100), .D(_1237__7_), .Q(Hhash_synth1_7_) );
	DFFPOSX1 DFFPOSX1_927 ( .CLK(clk_bF_buf99), .D(_1237__8_), .Q(Hhash_synth1_8_) );
	DFFPOSX1 DFFPOSX1_928 ( .CLK(clk_bF_buf98), .D(_1237__9_), .Q(Hhash_synth1_9_) );
	DFFPOSX1 DFFPOSX1_929 ( .CLK(clk_bF_buf97), .D(_1237__10_), .Q(Hhash_synth1_10_) );
	DFFPOSX1 DFFPOSX1_930 ( .CLK(clk_bF_buf96), .D(_1237__11_), .Q(Hhash_synth1_11_) );
	DFFPOSX1 DFFPOSX1_931 ( .CLK(clk_bF_buf95), .D(_1237__12_), .Q(Hhash_synth1_12_) );
	DFFPOSX1 DFFPOSX1_932 ( .CLK(clk_bF_buf94), .D(_1237__13_), .Q(Hhash_synth1_13_) );
	DFFPOSX1 DFFPOSX1_933 ( .CLK(clk_bF_buf93), .D(_1237__14_), .Q(Hhash_synth1_14_) );
	DFFPOSX1 DFFPOSX1_934 ( .CLK(clk_bF_buf92), .D(_1237__15_), .Q(Hhash_synth1_15_) );
	DFFPOSX1 DFFPOSX1_935 ( .CLK(clk_bF_buf91), .D(_1237__16_), .Q(Hhash_synth1_16_) );
	DFFPOSX1 DFFPOSX1_936 ( .CLK(clk_bF_buf90), .D(_1237__17_), .Q(Hhash_synth1_17_) );
	DFFPOSX1 DFFPOSX1_937 ( .CLK(clk_bF_buf89), .D(_1237__18_), .Q(Hhash_synth1_18_) );
	DFFPOSX1 DFFPOSX1_938 ( .CLK(clk_bF_buf88), .D(_1237__19_), .Q(Hhash_synth1_19_) );
	DFFPOSX1 DFFPOSX1_939 ( .CLK(clk_bF_buf87), .D(_1237__20_), .Q(Hhash_synth1_20_) );
	DFFPOSX1 DFFPOSX1_940 ( .CLK(clk_bF_buf86), .D(_1237__21_), .Q(Hhash_synth1_21_) );
	DFFPOSX1 DFFPOSX1_941 ( .CLK(clk_bF_buf85), .D(_1237__22_), .Q(Hhash_synth1_22_) );
	DFFPOSX1 DFFPOSX1_942 ( .CLK(clk_bF_buf84), .D(_1237__23_), .Q(Hhash_synth1_23_) );
	DFFPOSX1 DFFPOSX1_943 ( .CLK(clk_bF_buf83), .D(_1242__0_), .Q(micro_hash_synth_1_nonce_synth_1_0_) );
	DFFPOSX1 DFFPOSX1_944 ( .CLK(clk_bF_buf82), .D(_1242__1_), .Q(micro_hash_synth_1_nonce_synth_1_1_) );
	DFFPOSX1 DFFPOSX1_945 ( .CLK(clk_bF_buf81), .D(_1242__2_), .Q(micro_hash_synth_1_nonce_synth_1_2_) );
	DFFPOSX1 DFFPOSX1_946 ( .CLK(clk_bF_buf80), .D(_1242__3_), .Q(micro_hash_synth_1_nonce_synth_1_3_) );
	DFFPOSX1 DFFPOSX1_947 ( .CLK(clk_bF_buf79), .D(_1242__4_), .Q(micro_hash_synth_1_nonce_synth_1_4_) );
	DFFPOSX1 DFFPOSX1_948 ( .CLK(clk_bF_buf78), .D(_1242__5_), .Q(micro_hash_synth_1_nonce_synth_1_5_) );
	DFFPOSX1 DFFPOSX1_949 ( .CLK(clk_bF_buf77), .D(_1242__6_), .Q(micro_hash_synth_1_nonce_synth_1_6_) );
	DFFPOSX1 DFFPOSX1_950 ( .CLK(clk_bF_buf76), .D(_1242__7_), .Q(micro_hash_synth_1_nonce_synth_1_7_) );
	DFFPOSX1 DFFPOSX1_951 ( .CLK(clk_bF_buf75), .D(_1242__8_), .Q(micro_hash_synth_1_nonce_synth_1_8_) );
	DFFPOSX1 DFFPOSX1_952 ( .CLK(clk_bF_buf74), .D(_1242__9_), .Q(micro_hash_synth_1_nonce_synth_1_9_) );
	DFFPOSX1 DFFPOSX1_953 ( .CLK(clk_bF_buf73), .D(_1242__10_), .Q(micro_hash_synth_1_nonce_synth_1_10_) );
	DFFPOSX1 DFFPOSX1_954 ( .CLK(clk_bF_buf72), .D(_1242__11_), .Q(micro_hash_synth_1_nonce_synth_1_11_) );
	DFFPOSX1 DFFPOSX1_955 ( .CLK(clk_bF_buf71), .D(_1242__12_), .Q(micro_hash_synth_1_nonce_synth_1_12_) );
	DFFPOSX1 DFFPOSX1_956 ( .CLK(clk_bF_buf70), .D(_1242__13_), .Q(micro_hash_synth_1_nonce_synth_1_13_) );
	DFFPOSX1 DFFPOSX1_957 ( .CLK(clk_bF_buf69), .D(_1242__14_), .Q(micro_hash_synth_1_nonce_synth_1_14_) );
	DFFPOSX1 DFFPOSX1_958 ( .CLK(clk_bF_buf68), .D(_1242__15_), .Q(micro_hash_synth_1_nonce_synth_1_15_) );
	DFFPOSX1 DFFPOSX1_959 ( .CLK(clk_bF_buf67), .D(_1242__16_), .Q(micro_hash_synth_1_nonce_synth_1_16_) );
	DFFPOSX1 DFFPOSX1_960 ( .CLK(clk_bF_buf66), .D(_1242__17_), .Q(micro_hash_synth_1_nonce_synth_1_17_) );
	DFFPOSX1 DFFPOSX1_961 ( .CLK(clk_bF_buf65), .D(_1242__18_), .Q(micro_hash_synth_1_nonce_synth_1_18_) );
	DFFPOSX1 DFFPOSX1_962 ( .CLK(clk_bF_buf64), .D(_1242__19_), .Q(micro_hash_synth_1_nonce_synth_1_19_) );
	DFFPOSX1 DFFPOSX1_963 ( .CLK(clk_bF_buf63), .D(_1242__20_), .Q(micro_hash_synth_1_nonce_synth_1_20_) );
	DFFPOSX1 DFFPOSX1_964 ( .CLK(clk_bF_buf62), .D(_1242__21_), .Q(micro_hash_synth_1_nonce_synth_1_21_) );
	DFFPOSX1 DFFPOSX1_965 ( .CLK(clk_bF_buf61), .D(_1242__22_), .Q(micro_hash_synth_1_nonce_synth_1_22_) );
	DFFPOSX1 DFFPOSX1_966 ( .CLK(clk_bF_buf60), .D(_1242__23_), .Q(micro_hash_synth_1_nonce_synth_1_23_) );
	DFFPOSX1 DFFPOSX1_967 ( .CLK(clk_bF_buf59), .D(_1242__24_), .Q(micro_hash_synth_1_nonce_synth_1_24_) );
	DFFPOSX1 DFFPOSX1_968 ( .CLK(clk_bF_buf58), .D(_1242__25_), .Q(micro_hash_synth_1_nonce_synth_1_25_) );
	DFFPOSX1 DFFPOSX1_969 ( .CLK(clk_bF_buf57), .D(_1242__26_), .Q(micro_hash_synth_1_nonce_synth_1_26_) );
	DFFPOSX1 DFFPOSX1_970 ( .CLK(clk_bF_buf56), .D(_1242__27_), .Q(micro_hash_synth_1_nonce_synth_1_27_) );
	DFFPOSX1 DFFPOSX1_971 ( .CLK(clk_bF_buf55), .D(_1242__28_), .Q(micro_hash_synth_1_nonce_synth_1_28_) );
	DFFPOSX1 DFFPOSX1_972 ( .CLK(clk_bF_buf54), .D(_1242__29_), .Q(micro_hash_synth_1_nonce_synth_1_29_) );
	DFFPOSX1 DFFPOSX1_973 ( .CLK(clk_bF_buf53), .D(_1242__30_), .Q(micro_hash_synth_1_nonce_synth_1_30_) );
	DFFPOSX1 DFFPOSX1_974 ( .CLK(clk_bF_buf52), .D(_1242__31_), .Q(micro_hash_synth_1_nonce_synth_1_31_) );
	DFFPOSX1 DFFPOSX1_975 ( .CLK(clk_bF_buf51), .D(_1238__0_), .Q(micro_hash_synth_1_a_0_) );
	DFFPOSX1 DFFPOSX1_976 ( .CLK(clk_bF_buf50), .D(_1238__1_), .Q(micro_hash_synth_1_a_1_) );
	DFFPOSX1 DFFPOSX1_977 ( .CLK(clk_bF_buf49), .D(_1238__2_), .Q(micro_hash_synth_1_a_2_) );
	DFFPOSX1 DFFPOSX1_978 ( .CLK(clk_bF_buf48), .D(_1238__3_), .Q(micro_hash_synth_1_a_3_) );
	DFFPOSX1 DFFPOSX1_979 ( .CLK(clk_bF_buf47), .D(_1238__4_), .Q(micro_hash_synth_1_a_4_) );
	DFFPOSX1 DFFPOSX1_980 ( .CLK(clk_bF_buf46), .D(_1238__5_), .Q(micro_hash_synth_1_a_5_) );
	DFFPOSX1 DFFPOSX1_981 ( .CLK(clk_bF_buf45), .D(_1238__6_), .Q(micro_hash_synth_1_a_6_) );
	DFFPOSX1 DFFPOSX1_982 ( .CLK(clk_bF_buf44), .D(_1238__7_), .Q(micro_hash_synth_1_a_7_) );
	DFFPOSX1 DFFPOSX1_983 ( .CLK(clk_bF_buf43), .D(_1239__0_), .Q(micro_hash_synth_1_b_0_) );
	DFFPOSX1 DFFPOSX1_984 ( .CLK(clk_bF_buf42), .D(_1239__1_), .Q(micro_hash_synth_1_b_1_) );
	DFFPOSX1 DFFPOSX1_985 ( .CLK(clk_bF_buf41), .D(_1239__2_), .Q(micro_hash_synth_1_b_2_) );
	DFFPOSX1 DFFPOSX1_986 ( .CLK(clk_bF_buf40), .D(_1239__3_), .Q(micro_hash_synth_1_b_3_) );
	DFFPOSX1 DFFPOSX1_987 ( .CLK(clk_bF_buf39), .D(_1239__4_), .Q(micro_hash_synth_1_b_4_) );
	DFFPOSX1 DFFPOSX1_988 ( .CLK(clk_bF_buf38), .D(_1239__5_), .Q(micro_hash_synth_1_b_5_) );
	DFFPOSX1 DFFPOSX1_989 ( .CLK(clk_bF_buf37), .D(_1239__6_), .Q(micro_hash_synth_1_b_6_) );
	DFFPOSX1 DFFPOSX1_990 ( .CLK(clk_bF_buf36), .D(_1239__7_), .Q(micro_hash_synth_1_b_7_) );
	DFFPOSX1 DFFPOSX1_991 ( .CLK(clk_bF_buf35), .D(_1240__0_), .Q(micro_hash_synth_1_c_0_) );
	DFFPOSX1 DFFPOSX1_992 ( .CLK(clk_bF_buf34), .D(_1240__1_), .Q(micro_hash_synth_1_c_1_) );
	DFFPOSX1 DFFPOSX1_993 ( .CLK(clk_bF_buf33), .D(_1240__2_), .Q(micro_hash_synth_1_c_2_) );
	DFFPOSX1 DFFPOSX1_994 ( .CLK(clk_bF_buf32), .D(_1240__3_), .Q(micro_hash_synth_1_c_3_) );
	DFFPOSX1 DFFPOSX1_995 ( .CLK(clk_bF_buf31), .D(_1240__4_), .Q(micro_hash_synth_1_c_4_) );
	DFFPOSX1 DFFPOSX1_996 ( .CLK(clk_bF_buf30), .D(_1240__5_), .Q(micro_hash_synth_1_c_5_) );
	DFFPOSX1 DFFPOSX1_997 ( .CLK(clk_bF_buf29), .D(_1240__6_), .Q(micro_hash_synth_1_c_6_) );
	DFFPOSX1 DFFPOSX1_998 ( .CLK(clk_bF_buf28), .D(_1240__7_), .Q(micro_hash_synth_1_c_7_) );
	DFFPOSX1 DFFPOSX1_999 ( .CLK(clk_bF_buf27), .D(_1241__0_), .Q(micro_hash_synth_1_k_0_) );
	DFFPOSX1 DFFPOSX1_1000 ( .CLK(clk_bF_buf26), .D(_1241__1_), .Q(micro_hash_synth_1_k_1_) );
	DFFPOSX1 DFFPOSX1_1001 ( .CLK(clk_bF_buf25), .D(_1241__2_), .Q(micro_hash_synth_1_k_2_) );
	DFFPOSX1 DFFPOSX1_1002 ( .CLK(clk_bF_buf24), .D(_1241__3_), .Q(micro_hash_synth_1_k_3_) );
	DFFPOSX1 DFFPOSX1_1003 ( .CLK(clk_bF_buf23), .D(_1241__4_), .Q(micro_hash_synth_1_k_4_) );
	DFFPOSX1 DFFPOSX1_1004 ( .CLK(clk_bF_buf22), .D(_1241__5_), .Q(micro_hash_synth_1_k_5_) );
	DFFPOSX1 DFFPOSX1_1005 ( .CLK(clk_bF_buf21), .D(_1241__6_), .Q(micro_hash_synth_1_k_6_) );
	DFFPOSX1 DFFPOSX1_1006 ( .CLK(clk_bF_buf20), .D(_1241__7_), .Q(micro_hash_synth_1_k_7_) );
	DFFPOSX1 DFFPOSX1_1007 ( .CLK(clk_bF_buf19), .D(_1243__0_), .Q(micro_hash_synth_1_x_0_) );
	DFFPOSX1 DFFPOSX1_1008 ( .CLK(clk_bF_buf18), .D(_1243__1_), .Q(micro_hash_synth_1_x_1_) );
	DFFPOSX1 DFFPOSX1_1009 ( .CLK(clk_bF_buf17), .D(_1243__2_), .Q(micro_hash_synth_1_x_2_) );
	DFFPOSX1 DFFPOSX1_1010 ( .CLK(clk_bF_buf16), .D(_1243__3_), .Q(micro_hash_synth_1_x_3_) );
	DFFPOSX1 DFFPOSX1_1011 ( .CLK(clk_bF_buf15), .D(_1243__4_), .Q(micro_hash_synth_1_x_4_) );
	DFFPOSX1 DFFPOSX1_1012 ( .CLK(clk_bF_buf14), .D(_1243__5_), .Q(micro_hash_synth_1_x_5_) );
	DFFPOSX1 DFFPOSX1_1013 ( .CLK(clk_bF_buf13), .D(_1243__6_), .Q(micro_hash_synth_1_x_6_) );
	DFFPOSX1 DFFPOSX1_1014 ( .CLK(clk_bF_buf12), .D(_1243__7_), .Q(micro_hash_synth_1_x_7_) );
	DFFPOSX1 DFFPOSX1_1015 ( .CLK(clk_bF_buf11), .D(_1276_), .Q(micro_hash_synth_1_W_18__0_) );
	DFFPOSX1 DFFPOSX1_1016 ( .CLK(clk_bF_buf10), .D(_1277_), .Q(micro_hash_synth_1_W_18__1_) );
	DFFPOSX1 DFFPOSX1_1017 ( .CLK(clk_bF_buf9), .D(_1278_), .Q(micro_hash_synth_1_W_18__2_) );
	DFFPOSX1 DFFPOSX1_1018 ( .CLK(clk_bF_buf8), .D(_1279_), .Q(micro_hash_synth_1_W_18__3_) );
	DFFPOSX1 DFFPOSX1_1019 ( .CLK(clk_bF_buf7), .D(_1280_), .Q(micro_hash_synth_1_W_18__4_) );
	DFFPOSX1 DFFPOSX1_1020 ( .CLK(clk_bF_buf6), .D(_1281_), .Q(micro_hash_synth_1_W_18__5_) );
	DFFPOSX1 DFFPOSX1_1021 ( .CLK(clk_bF_buf5), .D(_1282_), .Q(micro_hash_synth_1_W_18__6_) );
	DFFPOSX1 DFFPOSX1_1022 ( .CLK(clk_bF_buf4), .D(_1283_), .Q(micro_hash_synth_1_W_18__7_) );
	DFFPOSX1 DFFPOSX1_1023 ( .CLK(clk_bF_buf3), .D(_1284_), .Q(micro_hash_synth_1_W_17__0_) );
	DFFPOSX1 DFFPOSX1_1024 ( .CLK(clk_bF_buf2), .D(_1286_), .Q(micro_hash_synth_1_W_17__1_) );
	DFFPOSX1 DFFPOSX1_1025 ( .CLK(clk_bF_buf1), .D(_1287_), .Q(micro_hash_synth_1_W_17__2_) );
	DFFPOSX1 DFFPOSX1_1026 ( .CLK(clk_bF_buf0), .D(_1288_), .Q(micro_hash_synth_1_W_17__3_) );
	DFFPOSX1 DFFPOSX1_1027 ( .CLK(clk_bF_buf113), .D(_1289_), .Q(micro_hash_synth_1_W_17__4_) );
	DFFPOSX1 DFFPOSX1_1028 ( .CLK(clk_bF_buf112), .D(_1290_), .Q(micro_hash_synth_1_W_17__5_) );
	DFFPOSX1 DFFPOSX1_1029 ( .CLK(clk_bF_buf111), .D(_1291_), .Q(micro_hash_synth_1_W_17__6_) );
	DFFPOSX1 DFFPOSX1_1030 ( .CLK(clk_bF_buf110), .D(_1292_), .Q(micro_hash_synth_1_W_17__7_) );
	DFFPOSX1 DFFPOSX1_1031 ( .CLK(clk_bF_buf109), .D(_1319_), .Q(micro_hash_synth_1_W_16__0_) );
	DFFPOSX1 DFFPOSX1_1032 ( .CLK(clk_bF_buf108), .D(_1320_), .Q(micro_hash_synth_1_W_16__1_) );
	DFFPOSX1 DFFPOSX1_1033 ( .CLK(clk_bF_buf107), .D(_1321_), .Q(micro_hash_synth_1_W_16__2_) );
	DFFPOSX1 DFFPOSX1_1034 ( .CLK(clk_bF_buf106), .D(_1322_), .Q(micro_hash_synth_1_W_16__3_) );
	DFFPOSX1 DFFPOSX1_1035 ( .CLK(clk_bF_buf105), .D(_1323_), .Q(micro_hash_synth_1_W_16__4_) );
	DFFPOSX1 DFFPOSX1_1036 ( .CLK(clk_bF_buf104), .D(_1324_), .Q(micro_hash_synth_1_W_16__5_) );
	DFFPOSX1 DFFPOSX1_1037 ( .CLK(clk_bF_buf103), .D(_1325_), .Q(micro_hash_synth_1_W_16__6_) );
	DFFPOSX1 DFFPOSX1_1038 ( .CLK(clk_bF_buf102), .D(_1326_), .Q(micro_hash_synth_1_W_16__7_) );
	DFFPOSX1 DFFPOSX1_1039 ( .CLK(clk_bF_buf101), .D(_1293_), .Q(micro_hash_synth_1_W_15__0_) );
	DFFPOSX1 DFFPOSX1_1040 ( .CLK(clk_bF_buf100), .D(_1294_), .Q(micro_hash_synth_1_W_15__1_) );
	DFFPOSX1 DFFPOSX1_1041 ( .CLK(clk_bF_buf99), .D(_1295_), .Q(micro_hash_synth_1_W_15__2_) );
	DFFPOSX1 DFFPOSX1_1042 ( .CLK(clk_bF_buf98), .D(_1296_), .Q(micro_hash_synth_1_W_15__3_) );
	DFFPOSX1 DFFPOSX1_1043 ( .CLK(clk_bF_buf97), .D(_1297_), .Q(micro_hash_synth_1_W_15__4_) );
	DFFPOSX1 DFFPOSX1_1044 ( .CLK(clk_bF_buf96), .D(_1298_), .Q(micro_hash_synth_1_W_15__5_) );
	DFFPOSX1 DFFPOSX1_1045 ( .CLK(clk_bF_buf95), .D(_1299_), .Q(micro_hash_synth_1_W_15__6_) );
	DFFPOSX1 DFFPOSX1_1046 ( .CLK(clk_bF_buf94), .D(_1300_), .Q(micro_hash_synth_1_W_15__7_) );
	DFFPOSX1 DFFPOSX1_1047 ( .CLK(clk_bF_buf93), .D(_1258_), .Q(micro_hash_synth_1_W_14__0_) );
	DFFPOSX1 DFFPOSX1_1048 ( .CLK(clk_bF_buf92), .D(_1259_), .Q(micro_hash_synth_1_W_14__1_) );
	DFFPOSX1 DFFPOSX1_1049 ( .CLK(clk_bF_buf91), .D(_1260_), .Q(micro_hash_synth_1_W_14__2_) );
	DFFPOSX1 DFFPOSX1_1050 ( .CLK(clk_bF_buf90), .D(_1261_), .Q(micro_hash_synth_1_W_14__3_) );
	DFFPOSX1 DFFPOSX1_1051 ( .CLK(clk_bF_buf89), .D(_1262_), .Q(micro_hash_synth_1_W_14__4_) );
	DFFPOSX1 DFFPOSX1_1052 ( .CLK(clk_bF_buf88), .D(_1263_), .Q(micro_hash_synth_1_W_14__5_) );
	DFFPOSX1 DFFPOSX1_1053 ( .CLK(clk_bF_buf87), .D(_1264_), .Q(micro_hash_synth_1_W_14__6_) );
	DFFPOSX1 DFFPOSX1_1054 ( .CLK(clk_bF_buf86), .D(_1265_), .Q(micro_hash_synth_1_W_14__7_) );
	DFFPOSX1 DFFPOSX1_1055 ( .CLK(clk_bF_buf85), .D(_1310_), .Q(micro_hash_synth_1_W_13__0_) );
	DFFPOSX1 DFFPOSX1_1056 ( .CLK(clk_bF_buf84), .D(_1311_), .Q(micro_hash_synth_1_W_13__1_) );
	DFFPOSX1 DFFPOSX1_1057 ( .CLK(clk_bF_buf83), .D(_1312_), .Q(micro_hash_synth_1_W_13__2_) );
	DFFPOSX1 DFFPOSX1_1058 ( .CLK(clk_bF_buf82), .D(_1313_), .Q(micro_hash_synth_1_W_13__3_) );
	DFFPOSX1 DFFPOSX1_1059 ( .CLK(clk_bF_buf81), .D(_1314_), .Q(micro_hash_synth_1_W_13__4_) );
	DFFPOSX1 DFFPOSX1_1060 ( .CLK(clk_bF_buf80), .D(_1315_), .Q(micro_hash_synth_1_W_13__5_) );
	DFFPOSX1 DFFPOSX1_1061 ( .CLK(clk_bF_buf79), .D(_1316_), .Q(micro_hash_synth_1_W_13__6_) );
	DFFPOSX1 DFFPOSX1_1062 ( .CLK(clk_bF_buf78), .D(_1318_), .Q(micro_hash_synth_1_W_13__7_) );
	DFFPOSX1 DFFPOSX1_1063 ( .CLK(clk_bF_buf77), .D(_1476_), .Q(micro_hash_synth_1_W_12__0_) );
	DFFPOSX1 DFFPOSX1_1064 ( .CLK(clk_bF_buf76), .D(_1477_), .Q(micro_hash_synth_1_W_12__1_) );
	DFFPOSX1 DFFPOSX1_1065 ( .CLK(clk_bF_buf75), .D(_1479_), .Q(micro_hash_synth_1_W_12__2_) );
	DFFPOSX1 DFFPOSX1_1066 ( .CLK(clk_bF_buf74), .D(_1480_), .Q(micro_hash_synth_1_W_12__3_) );
	DFFPOSX1 DFFPOSX1_1067 ( .CLK(clk_bF_buf73), .D(_1481_), .Q(micro_hash_synth_1_W_12__4_) );
	DFFPOSX1 DFFPOSX1_1068 ( .CLK(clk_bF_buf72), .D(_1482_), .Q(micro_hash_synth_1_W_12__5_) );
	DFFPOSX1 DFFPOSX1_1069 ( .CLK(clk_bF_buf71), .D(_1483_), .Q(micro_hash_synth_1_W_12__6_) );
	DFFPOSX1 DFFPOSX1_1070 ( .CLK(clk_bF_buf70), .D(_1484_), .Q(micro_hash_synth_1_W_12__7_) );
	DFFPOSX1 DFFPOSX1_1071 ( .CLK(clk_bF_buf69), .D(_1344_), .Q(micro_hash_synth_1_W_11__0_) );
	DFFPOSX1 DFFPOSX1_1072 ( .CLK(clk_bF_buf68), .D(_1345_), .Q(micro_hash_synth_1_W_11__1_) );
	DFFPOSX1 DFFPOSX1_1073 ( .CLK(clk_bF_buf67), .D(_1346_), .Q(micro_hash_synth_1_W_11__2_) );
	DFFPOSX1 DFFPOSX1_1074 ( .CLK(clk_bF_buf66), .D(_1347_), .Q(micro_hash_synth_1_W_11__3_) );
	DFFPOSX1 DFFPOSX1_1075 ( .CLK(clk_bF_buf65), .D(_1348_), .Q(micro_hash_synth_1_W_11__4_) );
	DFFPOSX1 DFFPOSX1_1076 ( .CLK(clk_bF_buf64), .D(_1349_), .Q(micro_hash_synth_1_W_11__5_) );
	DFFPOSX1 DFFPOSX1_1077 ( .CLK(clk_bF_buf63), .D(_1350_), .Q(micro_hash_synth_1_W_11__6_) );
	DFFPOSX1 DFFPOSX1_1078 ( .CLK(clk_bF_buf62), .D(_1351_), .Q(micro_hash_synth_1_W_11__7_) );
	DFFPOSX1 DFFPOSX1_1079 ( .CLK(clk_bF_buf61), .D(_1336_), .Q(micro_hash_synth_1_W_10__0_) );
	DFFPOSX1 DFFPOSX1_1080 ( .CLK(clk_bF_buf60), .D(_1337_), .Q(micro_hash_synth_1_W_10__1_) );
	DFFPOSX1 DFFPOSX1_1081 ( .CLK(clk_bF_buf59), .D(_1338_), .Q(micro_hash_synth_1_W_10__2_) );
	DFFPOSX1 DFFPOSX1_1082 ( .CLK(clk_bF_buf58), .D(_1339_), .Q(micro_hash_synth_1_W_10__3_) );
	DFFPOSX1 DFFPOSX1_1083 ( .CLK(clk_bF_buf57), .D(_1340_), .Q(micro_hash_synth_1_W_10__4_) );
	DFFPOSX1 DFFPOSX1_1084 ( .CLK(clk_bF_buf56), .D(_1341_), .Q(micro_hash_synth_1_W_10__5_) );
	DFFPOSX1 DFFPOSX1_1085 ( .CLK(clk_bF_buf55), .D(_1342_), .Q(micro_hash_synth_1_W_10__6_) );
	DFFPOSX1 DFFPOSX1_1086 ( .CLK(clk_bF_buf54), .D(_1343_), .Q(micro_hash_synth_1_W_10__7_) );
	DFFPOSX1 DFFPOSX1_1087 ( .CLK(clk_bF_buf53), .D(_1441_), .Q(micro_hash_synth_1_W_9__0_) );
	DFFPOSX1 DFFPOSX1_1088 ( .CLK(clk_bF_buf52), .D(_1442_), .Q(micro_hash_synth_1_W_9__1_) );
	DFFPOSX1 DFFPOSX1_1089 ( .CLK(clk_bF_buf51), .D(_1443_), .Q(micro_hash_synth_1_W_9__2_) );
	DFFPOSX1 DFFPOSX1_1090 ( .CLK(clk_bF_buf50), .D(_1444_), .Q(micro_hash_synth_1_W_9__3_) );
	DFFPOSX1 DFFPOSX1_1091 ( .CLK(clk_bF_buf49), .D(_1446_), .Q(micro_hash_synth_1_W_9__4_) );
	DFFPOSX1 DFFPOSX1_1092 ( .CLK(clk_bF_buf48), .D(_1447_), .Q(micro_hash_synth_1_W_9__5_) );
	DFFPOSX1 DFFPOSX1_1093 ( .CLK(clk_bF_buf47), .D(_1448_), .Q(micro_hash_synth_1_W_9__6_) );
	DFFPOSX1 DFFPOSX1_1094 ( .CLK(clk_bF_buf46), .D(_1449_), .Q(micro_hash_synth_1_W_9__7_) );
	DFFPOSX1 DFFPOSX1_1095 ( .CLK(clk_bF_buf45), .D(_1492_), .Q(micro_hash_synth_1_W_8__0_) );
	DFFPOSX1 DFFPOSX1_1096 ( .CLK(clk_bF_buf44), .D(_1497_), .Q(micro_hash_synth_1_W_8__1_) );
	DFFPOSX1 DFFPOSX1_1097 ( .CLK(clk_bF_buf43), .D(_1498_), .Q(micro_hash_synth_1_W_8__2_) );
	DFFPOSX1 DFFPOSX1_1098 ( .CLK(clk_bF_buf42), .D(_1499_), .Q(micro_hash_synth_1_W_8__3_) );
	DFFPOSX1 DFFPOSX1_1099 ( .CLK(clk_bF_buf41), .D(_1244_), .Q(micro_hash_synth_1_W_8__4_) );
	DFFPOSX1 DFFPOSX1_1100 ( .CLK(clk_bF_buf40), .D(_1245_), .Q(micro_hash_synth_1_W_8__5_) );
	DFFPOSX1 DFFPOSX1_1101 ( .CLK(clk_bF_buf39), .D(_1253_), .Q(micro_hash_synth_1_W_8__6_) );
	DFFPOSX1 DFFPOSX1_1102 ( .CLK(clk_bF_buf38), .D(_1255_), .Q(micro_hash_synth_1_W_8__7_) );
	DFFPOSX1 DFFPOSX1_1103 ( .CLK(clk_bF_buf37), .D(_1424_), .Q(micro_hash_synth_1_W_7__0_) );
	DFFPOSX1 DFFPOSX1_1104 ( .CLK(clk_bF_buf36), .D(_1425_), .Q(micro_hash_synth_1_W_7__1_) );
	DFFPOSX1 DFFPOSX1_1105 ( .CLK(clk_bF_buf35), .D(_1426_), .Q(micro_hash_synth_1_W_7__2_) );
	DFFPOSX1 DFFPOSX1_1106 ( .CLK(clk_bF_buf34), .D(_1427_), .Q(micro_hash_synth_1_W_7__3_) );
	DFFPOSX1 DFFPOSX1_1107 ( .CLK(clk_bF_buf33), .D(_1428_), .Q(micro_hash_synth_1_W_7__4_) );
	DFFPOSX1 DFFPOSX1_1108 ( .CLK(clk_bF_buf32), .D(_1429_), .Q(micro_hash_synth_1_W_7__5_) );
	DFFPOSX1 DFFPOSX1_1109 ( .CLK(clk_bF_buf31), .D(_1430_), .Q(micro_hash_synth_1_W_7__6_) );
	DFFPOSX1 DFFPOSX1_1110 ( .CLK(clk_bF_buf30), .D(_1431_), .Q(micro_hash_synth_1_W_7__7_) );
	DFFPOSX1 DFFPOSX1_1111 ( .CLK(clk_bF_buf29), .D(_1302_), .Q(micro_hash_synth_1_W_6__0_) );
	DFFPOSX1 DFFPOSX1_1112 ( .CLK(clk_bF_buf28), .D(_1303_), .Q(micro_hash_synth_1_W_6__1_) );
	DFFPOSX1 DFFPOSX1_1113 ( .CLK(clk_bF_buf27), .D(_1304_), .Q(micro_hash_synth_1_W_6__2_) );
	DFFPOSX1 DFFPOSX1_1114 ( .CLK(clk_bF_buf26), .D(_1305_), .Q(micro_hash_synth_1_W_6__3_) );
	DFFPOSX1 DFFPOSX1_1115 ( .CLK(clk_bF_buf25), .D(_1306_), .Q(micro_hash_synth_1_W_6__4_) );
	DFFPOSX1 DFFPOSX1_1116 ( .CLK(clk_bF_buf24), .D(_1307_), .Q(micro_hash_synth_1_W_6__5_) );
	DFFPOSX1 DFFPOSX1_1117 ( .CLK(clk_bF_buf23), .D(_1308_), .Q(micro_hash_synth_1_W_6__6_) );
	DFFPOSX1 DFFPOSX1_1118 ( .CLK(clk_bF_buf22), .D(_1309_), .Q(micro_hash_synth_1_W_6__7_) );
	DFFPOSX1 DFFPOSX1_1119 ( .CLK(clk_bF_buf21), .D(_1246_), .Q(micro_hash_synth_1_W_5__0_) );
	DFFPOSX1 DFFPOSX1_1120 ( .CLK(clk_bF_buf20), .D(_1247_), .Q(micro_hash_synth_1_W_5__1_) );
	DFFPOSX1 DFFPOSX1_1121 ( .CLK(clk_bF_buf19), .D(_1248_), .Q(micro_hash_synth_1_W_5__2_) );
	DFFPOSX1 DFFPOSX1_1122 ( .CLK(clk_bF_buf18), .D(_1249_), .Q(micro_hash_synth_1_W_5__3_) );
	DFFPOSX1 DFFPOSX1_1123 ( .CLK(clk_bF_buf17), .D(_1250_), .Q(micro_hash_synth_1_W_5__4_) );
	DFFPOSX1 DFFPOSX1_1124 ( .CLK(clk_bF_buf16), .D(_1251_), .Q(micro_hash_synth_1_W_5__5_) );
	DFFPOSX1 DFFPOSX1_1125 ( .CLK(clk_bF_buf15), .D(_1252_), .Q(micro_hash_synth_1_W_5__6_) );
	DFFPOSX1 DFFPOSX1_1126 ( .CLK(clk_bF_buf14), .D(_1254_), .Q(micro_hash_synth_1_W_5__7_) );
	DFFPOSX1 DFFPOSX1_1127 ( .CLK(clk_bF_buf13), .D(_1450_), .Q(micro_hash_synth_1_W_4__0_) );
	DFFPOSX1 DFFPOSX1_1128 ( .CLK(clk_bF_buf12), .D(_1451_), .Q(micro_hash_synth_1_W_4__1_) );
	DFFPOSX1 DFFPOSX1_1129 ( .CLK(clk_bF_buf11), .D(_1452_), .Q(micro_hash_synth_1_W_4__2_) );
	DFFPOSX1 DFFPOSX1_1130 ( .CLK(clk_bF_buf10), .D(_1453_), .Q(micro_hash_synth_1_W_4__3_) );
	DFFPOSX1 DFFPOSX1_1131 ( .CLK(clk_bF_buf9), .D(_1454_), .Q(micro_hash_synth_1_W_4__4_) );
	DFFPOSX1 DFFPOSX1_1132 ( .CLK(clk_bF_buf8), .D(_1455_), .Q(micro_hash_synth_1_W_4__5_) );
	DFFPOSX1 DFFPOSX1_1133 ( .CLK(clk_bF_buf7), .D(_1457_), .Q(micro_hash_synth_1_W_4__6_) );
	DFFPOSX1 DFFPOSX1_1134 ( .CLK(clk_bF_buf6), .D(_1458_), .Q(micro_hash_synth_1_W_4__7_) );
	DFFPOSX1 DFFPOSX1_1135 ( .CLK(clk_bF_buf5), .D(_1415_), .Q(micro_hash_synth_1_W_23__0_) );
	DFFPOSX1 DFFPOSX1_1136 ( .CLK(clk_bF_buf4), .D(_1416_), .Q(micro_hash_synth_1_W_23__1_) );
	DFFPOSX1 DFFPOSX1_1137 ( .CLK(clk_bF_buf3), .D(_1417_), .Q(micro_hash_synth_1_W_23__2_) );
	DFFPOSX1 DFFPOSX1_1138 ( .CLK(clk_bF_buf2), .D(_1418_), .Q(micro_hash_synth_1_W_23__3_) );
	DFFPOSX1 DFFPOSX1_1139 ( .CLK(clk_bF_buf1), .D(_1419_), .Q(micro_hash_synth_1_W_23__4_) );
	DFFPOSX1 DFFPOSX1_1140 ( .CLK(clk_bF_buf0), .D(_1420_), .Q(micro_hash_synth_1_W_23__5_) );
	DFFPOSX1 DFFPOSX1_1141 ( .CLK(clk_bF_buf113), .D(_1421_), .Q(micro_hash_synth_1_W_23__6_) );
	DFFPOSX1 DFFPOSX1_1142 ( .CLK(clk_bF_buf112), .D(_1422_), .Q(micro_hash_synth_1_W_23__7_) );
	DFFPOSX1 DFFPOSX1_1143 ( .CLK(clk_bF_buf111), .D(_1406_), .Q(micro_hash_synth_1_W_24__0_) );
	DFFPOSX1 DFFPOSX1_1144 ( .CLK(clk_bF_buf110), .D(_1407_), .Q(micro_hash_synth_1_W_24__1_) );
	DFFPOSX1 DFFPOSX1_1145 ( .CLK(clk_bF_buf109), .D(_1408_), .Q(micro_hash_synth_1_W_24__2_) );
	DFFPOSX1 DFFPOSX1_1146 ( .CLK(clk_bF_buf108), .D(_1409_), .Q(micro_hash_synth_1_W_24__3_) );
	DFFPOSX1 DFFPOSX1_1147 ( .CLK(clk_bF_buf107), .D(_1410_), .Q(micro_hash_synth_1_W_24__4_) );
	DFFPOSX1 DFFPOSX1_1148 ( .CLK(clk_bF_buf106), .D(_1411_), .Q(micro_hash_synth_1_W_24__5_) );
	DFFPOSX1 DFFPOSX1_1149 ( .CLK(clk_bF_buf105), .D(_1413_), .Q(micro_hash_synth_1_W_24__6_) );
	DFFPOSX1 DFFPOSX1_1150 ( .CLK(clk_bF_buf104), .D(_1414_), .Q(micro_hash_synth_1_W_24__7_) );
	DFFPOSX1 DFFPOSX1_1151 ( .CLK(clk_bF_buf103), .D(_1434_), .Q(micro_hash_synth_1_W_25__0_) );
	DFFPOSX1 DFFPOSX1_1152 ( .CLK(clk_bF_buf102), .D(_1445_), .Q(micro_hash_synth_1_W_25__1_) );
	DFFPOSX1 DFFPOSX1_1153 ( .CLK(clk_bF_buf101), .D(_1456_), .Q(micro_hash_synth_1_W_25__2_) );
	DFFPOSX1 DFFPOSX1_1154 ( .CLK(clk_bF_buf100), .D(_1467_), .Q(micro_hash_synth_1_W_25__3_) );
	DFFPOSX1 DFFPOSX1_1155 ( .CLK(clk_bF_buf99), .D(_1478_), .Q(micro_hash_synth_1_W_25__4_) );
	DFFPOSX1 DFFPOSX1_1156 ( .CLK(clk_bF_buf98), .D(_1485_), .Q(micro_hash_synth_1_W_25__5_) );
	DFFPOSX1 DFFPOSX1_1157 ( .CLK(clk_bF_buf97), .D(_1486_), .Q(micro_hash_synth_1_W_25__6_) );
	DFFPOSX1 DFFPOSX1_1158 ( .CLK(clk_bF_buf96), .D(_1487_), .Q(micro_hash_synth_1_W_25__7_) );
	DFFPOSX1 DFFPOSX1_1159 ( .CLK(clk_bF_buf95), .D(_1400_), .Q(micro_hash_synth_1_W_26__0_) );
	DFFPOSX1 DFFPOSX1_1160 ( .CLK(clk_bF_buf94), .D(_1401_), .Q(micro_hash_synth_1_W_26__1_) );
	DFFPOSX1 DFFPOSX1_1161 ( .CLK(clk_bF_buf93), .D(_1402_), .Q(micro_hash_synth_1_W_26__2_) );
	DFFPOSX1 DFFPOSX1_1162 ( .CLK(clk_bF_buf92), .D(_1403_), .Q(micro_hash_synth_1_W_26__3_) );
	DFFPOSX1 DFFPOSX1_1163 ( .CLK(clk_bF_buf91), .D(_1404_), .Q(micro_hash_synth_1_W_26__4_) );
	DFFPOSX1 DFFPOSX1_1164 ( .CLK(clk_bF_buf90), .D(_1405_), .Q(micro_hash_synth_1_W_26__5_) );
	DFFPOSX1 DFFPOSX1_1165 ( .CLK(clk_bF_buf89), .D(_1412_), .Q(micro_hash_synth_1_W_26__6_) );
	DFFPOSX1 DFFPOSX1_1166 ( .CLK(clk_bF_buf88), .D(_1423_), .Q(micro_hash_synth_1_W_26__7_) );
	DFFPOSX1 DFFPOSX1_1167 ( .CLK(clk_bF_buf87), .D(_1360_), .Q(micro_hash_synth_1_W_27__0_) );
	DFFPOSX1 DFFPOSX1_1168 ( .CLK(clk_bF_buf86), .D(_1361_), .Q(micro_hash_synth_1_W_27__1_) );
	DFFPOSX1 DFFPOSX1_1169 ( .CLK(clk_bF_buf85), .D(_1362_), .Q(micro_hash_synth_1_W_27__2_) );
	DFFPOSX1 DFFPOSX1_1170 ( .CLK(clk_bF_buf84), .D(_1363_), .Q(micro_hash_synth_1_W_27__3_) );
	DFFPOSX1 DFFPOSX1_1171 ( .CLK(clk_bF_buf83), .D(_1364_), .Q(micro_hash_synth_1_W_27__4_) );
	DFFPOSX1 DFFPOSX1_1172 ( .CLK(clk_bF_buf82), .D(_1365_), .Q(micro_hash_synth_1_W_27__5_) );
	DFFPOSX1 DFFPOSX1_1173 ( .CLK(clk_bF_buf81), .D(_1366_), .Q(micro_hash_synth_1_W_27__6_) );
	DFFPOSX1 DFFPOSX1_1174 ( .CLK(clk_bF_buf80), .D(_1367_), .Q(micro_hash_synth_1_W_27__7_) );
	DFFPOSX1 DFFPOSX1_1175 ( .CLK(clk_bF_buf79), .D(_1368_), .Q(micro_hash_synth_1_W_28__0_) );
	DFFPOSX1 DFFPOSX1_1176 ( .CLK(clk_bF_buf78), .D(_1369_), .Q(micro_hash_synth_1_W_28__1_) );
	DFFPOSX1 DFFPOSX1_1177 ( .CLK(clk_bF_buf77), .D(_1370_), .Q(micro_hash_synth_1_W_28__2_) );
	DFFPOSX1 DFFPOSX1_1178 ( .CLK(clk_bF_buf76), .D(_1371_), .Q(micro_hash_synth_1_W_28__3_) );
	DFFPOSX1 DFFPOSX1_1179 ( .CLK(clk_bF_buf75), .D(_1372_), .Q(micro_hash_synth_1_W_28__4_) );
	DFFPOSX1 DFFPOSX1_1180 ( .CLK(clk_bF_buf74), .D(_1373_), .Q(micro_hash_synth_1_W_28__5_) );
	DFFPOSX1 DFFPOSX1_1181 ( .CLK(clk_bF_buf73), .D(_1374_), .Q(micro_hash_synth_1_W_28__6_) );
	DFFPOSX1 DFFPOSX1_1182 ( .CLK(clk_bF_buf72), .D(_1375_), .Q(micro_hash_synth_1_W_28__7_) );
	DFFPOSX1 DFFPOSX1_1183 ( .CLK(clk_bF_buf71), .D(_1376_), .Q(micro_hash_synth_1_W_29__0_) );
	DFFPOSX1 DFFPOSX1_1184 ( .CLK(clk_bF_buf70), .D(_1377_), .Q(micro_hash_synth_1_W_29__1_) );
	DFFPOSX1 DFFPOSX1_1185 ( .CLK(clk_bF_buf69), .D(_1378_), .Q(micro_hash_synth_1_W_29__2_) );
	DFFPOSX1 DFFPOSX1_1186 ( .CLK(clk_bF_buf68), .D(_1379_), .Q(micro_hash_synth_1_W_29__3_) );
	DFFPOSX1 DFFPOSX1_1187 ( .CLK(clk_bF_buf67), .D(_1380_), .Q(micro_hash_synth_1_W_29__4_) );
	DFFPOSX1 DFFPOSX1_1188 ( .CLK(clk_bF_buf66), .D(_1381_), .Q(micro_hash_synth_1_W_29__5_) );
	DFFPOSX1 DFFPOSX1_1189 ( .CLK(clk_bF_buf65), .D(_1382_), .Q(micro_hash_synth_1_W_29__6_) );
	DFFPOSX1 DFFPOSX1_1190 ( .CLK(clk_bF_buf64), .D(_1383_), .Q(micro_hash_synth_1_W_29__7_) );
	DFFPOSX1 DFFPOSX1_1191 ( .CLK(clk_bF_buf63), .D(_1384_), .Q(micro_hash_synth_1_W_30__0_) );
	DFFPOSX1 DFFPOSX1_1192 ( .CLK(clk_bF_buf62), .D(_1385_), .Q(micro_hash_synth_1_W_30__1_) );
	DFFPOSX1 DFFPOSX1_1193 ( .CLK(clk_bF_buf61), .D(_1386_), .Q(micro_hash_synth_1_W_30__2_) );
	DFFPOSX1 DFFPOSX1_1194 ( .CLK(clk_bF_buf60), .D(_1387_), .Q(micro_hash_synth_1_W_30__3_) );
	DFFPOSX1 DFFPOSX1_1195 ( .CLK(clk_bF_buf59), .D(_1388_), .Q(micro_hash_synth_1_W_30__4_) );
	DFFPOSX1 DFFPOSX1_1196 ( .CLK(clk_bF_buf58), .D(_1389_), .Q(micro_hash_synth_1_W_30__5_) );
	DFFPOSX1 DFFPOSX1_1197 ( .CLK(clk_bF_buf57), .D(_1390_), .Q(micro_hash_synth_1_W_30__6_) );
	DFFPOSX1 DFFPOSX1_1198 ( .CLK(clk_bF_buf56), .D(_1391_), .Q(micro_hash_synth_1_W_30__7_) );
	DFFPOSX1 DFFPOSX1_1199 ( .CLK(clk_bF_buf55), .D(_1256_), .Q(micro_hash_synth_1_W_3__0_) );
	DFFPOSX1 DFFPOSX1_1200 ( .CLK(clk_bF_buf54), .D(_1257_), .Q(micro_hash_synth_1_W_3__1_) );
	DFFPOSX1 DFFPOSX1_1201 ( .CLK(clk_bF_buf53), .D(_1266_), .Q(micro_hash_synth_1_W_3__2_) );
	DFFPOSX1 DFFPOSX1_1202 ( .CLK(clk_bF_buf52), .D(_1269_), .Q(micro_hash_synth_1_W_3__3_) );
	DFFPOSX1 DFFPOSX1_1203 ( .CLK(clk_bF_buf51), .D(_1285_), .Q(micro_hash_synth_1_W_3__4_) );
	DFFPOSX1 DFFPOSX1_1204 ( .CLK(clk_bF_buf50), .D(_1301_), .Q(micro_hash_synth_1_W_3__5_) );
	DFFPOSX1 DFFPOSX1_1205 ( .CLK(clk_bF_buf49), .D(_1317_), .Q(micro_hash_synth_1_W_3__6_) );
	DFFPOSX1 DFFPOSX1_1206 ( .CLK(clk_bF_buf48), .D(_1333_), .Q(micro_hash_synth_1_W_3__7_) );
	DFFPOSX1 DFFPOSX1_1207 ( .CLK(clk_bF_buf47), .D(_1392_), .Q(micro_hash_synth_1_W_31__0_) );
	DFFPOSX1 DFFPOSX1_1208 ( .CLK(clk_bF_buf46), .D(_1393_), .Q(micro_hash_synth_1_W_31__1_) );
	DFFPOSX1 DFFPOSX1_1209 ( .CLK(clk_bF_buf45), .D(_1394_), .Q(micro_hash_synth_1_W_31__2_) );
	DFFPOSX1 DFFPOSX1_1210 ( .CLK(clk_bF_buf44), .D(_1395_), .Q(micro_hash_synth_1_W_31__3_) );
	DFFPOSX1 DFFPOSX1_1211 ( .CLK(clk_bF_buf43), .D(_1396_), .Q(micro_hash_synth_1_W_31__4_) );
	DFFPOSX1 DFFPOSX1_1212 ( .CLK(clk_bF_buf42), .D(_1397_), .Q(micro_hash_synth_1_W_31__5_) );
	DFFPOSX1 DFFPOSX1_1213 ( .CLK(clk_bF_buf41), .D(_1398_), .Q(micro_hash_synth_1_W_31__6_) );
	DFFPOSX1 DFFPOSX1_1214 ( .CLK(clk_bF_buf40), .D(_1399_), .Q(micro_hash_synth_1_W_31__7_) );
	DFFPOSX1 DFFPOSX1_1215 ( .CLK(clk_bF_buf39), .D(_1327_), .Q(micro_hash_synth_1_W_1__0_) );
	DFFPOSX1 DFFPOSX1_1216 ( .CLK(clk_bF_buf38), .D(_1328_), .Q(micro_hash_synth_1_W_1__1_) );
	DFFPOSX1 DFFPOSX1_1217 ( .CLK(clk_bF_buf37), .D(_1329_), .Q(micro_hash_synth_1_W_1__2_) );
	DFFPOSX1 DFFPOSX1_1218 ( .CLK(clk_bF_buf36), .D(_1330_), .Q(micro_hash_synth_1_W_1__3_) );
	DFFPOSX1 DFFPOSX1_1219 ( .CLK(clk_bF_buf35), .D(_1331_), .Q(micro_hash_synth_1_W_1__4_) );
	DFFPOSX1 DFFPOSX1_1220 ( .CLK(clk_bF_buf34), .D(_1332_), .Q(micro_hash_synth_1_W_1__5_) );
	DFFPOSX1 DFFPOSX1_1221 ( .CLK(clk_bF_buf33), .D(_1334_), .Q(micro_hash_synth_1_W_1__6_) );
	DFFPOSX1 DFFPOSX1_1222 ( .CLK(clk_bF_buf32), .D(_1335_), .Q(micro_hash_synth_1_W_1__7_) );
	DFFPOSX1 DFFPOSX1_1223 ( .CLK(clk_bF_buf31), .D(_1352_), .Q(micro_hash_synth_1_W_2__0_) );
	DFFPOSX1 DFFPOSX1_1224 ( .CLK(clk_bF_buf30), .D(_1353_), .Q(micro_hash_synth_1_W_2__1_) );
	DFFPOSX1 DFFPOSX1_1225 ( .CLK(clk_bF_buf29), .D(_1354_), .Q(micro_hash_synth_1_W_2__2_) );
	DFFPOSX1 DFFPOSX1_1226 ( .CLK(clk_bF_buf28), .D(_1355_), .Q(micro_hash_synth_1_W_2__3_) );
	DFFPOSX1 DFFPOSX1_1227 ( .CLK(clk_bF_buf27), .D(_1356_), .Q(micro_hash_synth_1_W_2__4_) );
	DFFPOSX1 DFFPOSX1_1228 ( .CLK(clk_bF_buf26), .D(_1357_), .Q(micro_hash_synth_1_W_2__5_) );
	DFFPOSX1 DFFPOSX1_1229 ( .CLK(clk_bF_buf25), .D(_1358_), .Q(micro_hash_synth_1_W_2__6_) );
	DFFPOSX1 DFFPOSX1_1230 ( .CLK(clk_bF_buf24), .D(_1359_), .Q(micro_hash_synth_1_W_2__7_) );
	INVX1 INVX1_1073 ( .A(micro_hash_synth_2_W_26__0_), .Y(_4728_) );
	OR2X2 OR2X2_57 ( .A(concatenador_counter_2d_3_), .B(concatenador_counter_2d_2_), .Y(_4729_) );
	NOR2X1 NOR2X1_473 ( .A(concatenador_counter_2d_5_), .B(concatenador_counter_2d_4_), .Y(_4730_) );
	INVX1 INVX1_1074 ( .A(_4730_), .Y(_4731_) );
	NOR2X1 NOR2X1_474 ( .A(_4729_), .B(_4731_), .Y(_4732_) );
	INVX8 INVX8_9 ( .A(concatenador_counter_2d_0_bF_buf7), .Y(_4733_) );
	NOR2X1 NOR2X1_475 ( .A(concatenador_counter_2d_1_bF_buf6), .B(_4733__bF_buf3), .Y(_4734_) );
	NAND3X1 NAND3X1_215 ( .A(reset_L_bF_buf0), .B(_4734_), .C(_4732_), .Y(_4735_) );
	NOR2X1 NOR2X1_476 ( .A(concatenador_counter_2d_1_bF_buf5), .B(_4729_), .Y(_4736_) );
	INVX1 INVX1_1075 ( .A(_4736_), .Y(_4737_) );
	NOR2X1 NOR2X1_477 ( .A(_4731_), .B(_4737_), .Y(_4738_) );
	INVX1 INVX1_1076 ( .A(_4738_), .Y(_4739_) );
	OAI21X1 OAI21X1_1218 ( .A(_4739_), .B(_4733__bF_buf2), .C(reset_L_bF_buf49), .Y(_4740_) );
	XOR2X1 XOR2X1_62 ( .A(micro_hash_synth_2_W_12__0_), .B(micro_hash_synth_2_W_17__0_), .Y(_4741_) );
	NOR2X1 NOR2X1_478 ( .A(micro_hash_synth_2_W_23__0_), .B(_4741_), .Y(_4742_) );
	OAI22X1 OAI22X1_477 ( .A(_4735__bF_buf15), .B(_4742_), .C(_4740__bF_buf12), .D(_4728_), .Y(_3210_) );
	INVX1 INVX1_1077 ( .A(micro_hash_synth_2_W_26__1_), .Y(_4743_) );
	INVX1 INVX1_1078 ( .A(micro_hash_synth_2_W_12__1_), .Y(_4744_) );
	INVX1 INVX1_1079 ( .A(micro_hash_synth_2_W_23__1_), .Y(_4745_) );
	OAI21X1 OAI21X1_1219 ( .A(_4744_), .B(micro_hash_synth_2_W_17__1_), .C(_4745_), .Y(_4746_) );
	AOI21X1 AOI21X1_850 ( .A(_4744_), .B(micro_hash_synth_2_W_17__1_), .C(_4746_), .Y(_4747_) );
	OAI22X1 OAI22X1_478 ( .A(_4735__bF_buf14), .B(_4747_), .C(_4740__bF_buf11), .D(_4743_), .Y(_3211_) );
	INVX1 INVX1_1080 ( .A(micro_hash_synth_2_W_26__2_), .Y(_4748_) );
	INVX1 INVX1_1081 ( .A(micro_hash_synth_2_W_12__2_), .Y(_4749_) );
	INVX1 INVX1_1082 ( .A(micro_hash_synth_2_W_23__2_), .Y(_4750_) );
	OAI21X1 OAI21X1_1220 ( .A(_4749_), .B(micro_hash_synth_2_W_17__2_), .C(_4750_), .Y(_4751_) );
	AOI21X1 AOI21X1_851 ( .A(_4749_), .B(micro_hash_synth_2_W_17__2_), .C(_4751_), .Y(_4752_) );
	OAI22X1 OAI22X1_479 ( .A(_4735__bF_buf13), .B(_4752_), .C(_4740__bF_buf10), .D(_4748_), .Y(_3212_) );
	INVX1 INVX1_1083 ( .A(micro_hash_synth_2_W_26__3_), .Y(_4753_) );
	XOR2X1 XOR2X1_63 ( .A(micro_hash_synth_2_W_12__3_), .B(micro_hash_synth_2_W_17__3_), .Y(_4754_) );
	NOR2X1 NOR2X1_479 ( .A(micro_hash_synth_2_W_23__3_), .B(_4754_), .Y(_4755_) );
	OAI22X1 OAI22X1_480 ( .A(_4735__bF_buf12), .B(_4755_), .C(_4740__bF_buf9), .D(_4753_), .Y(_3213_) );
	INVX1 INVX1_1084 ( .A(micro_hash_synth_2_W_26__4_), .Y(_4756_) );
	XOR2X1 XOR2X1_64 ( .A(micro_hash_synth_2_W_12__4_), .B(micro_hash_synth_2_W_17__4_), .Y(_4757_) );
	NOR2X1 NOR2X1_480 ( .A(micro_hash_synth_2_W_23__4_), .B(_4757_), .Y(_4758_) );
	OAI22X1 OAI22X1_481 ( .A(_4735__bF_buf11), .B(_4758_), .C(_4740__bF_buf8), .D(_4756_), .Y(_3214_) );
	INVX1 INVX1_1085 ( .A(micro_hash_synth_2_W_26__5_), .Y(_4759_) );
	XOR2X1 XOR2X1_65 ( .A(micro_hash_synth_2_W_12__5_), .B(micro_hash_synth_2_W_17__5_), .Y(_4760_) );
	NOR2X1 NOR2X1_481 ( .A(micro_hash_synth_2_W_23__5_), .B(_4760_), .Y(_4761_) );
	OAI22X1 OAI22X1_482 ( .A(_4735__bF_buf10), .B(_4761_), .C(_4740__bF_buf7), .D(_4759_), .Y(_3215_) );
	INVX1 INVX1_1086 ( .A(micro_hash_synth_2_W_26__6_), .Y(_4762_) );
	INVX1 INVX1_1087 ( .A(micro_hash_synth_2_W_12__6_), .Y(_4763_) );
	INVX1 INVX1_1088 ( .A(micro_hash_synth_2_W_23__6_), .Y(_4764_) );
	OAI21X1 OAI21X1_1221 ( .A(_4763_), .B(micro_hash_synth_2_W_17__6_), .C(_4764_), .Y(_4765_) );
	AOI21X1 AOI21X1_852 ( .A(_4763_), .B(micro_hash_synth_2_W_17__6_), .C(_4765_), .Y(_4766_) );
	OAI22X1 OAI22X1_483 ( .A(_4735__bF_buf9), .B(_4766_), .C(_4740__bF_buf6), .D(_4762_), .Y(_3222_) );
	INVX1 INVX1_1089 ( .A(micro_hash_synth_2_W_26__7_), .Y(_4767_) );
	INVX1 INVX1_1090 ( .A(micro_hash_synth_2_W_12__7_), .Y(_4768_) );
	INVX1 INVX1_1091 ( .A(micro_hash_synth_2_W_23__7_), .Y(_4769_) );
	OAI21X1 OAI21X1_1222 ( .A(_4768_), .B(micro_hash_synth_2_W_17__7_), .C(_4769_), .Y(_4770_) );
	AOI21X1 AOI21X1_853 ( .A(_4768_), .B(micro_hash_synth_2_W_17__7_), .C(_4770_), .Y(_4771_) );
	OAI22X1 OAI22X1_484 ( .A(_4735__bF_buf8), .B(_4771_), .C(_4740__bF_buf5), .D(_4767_), .Y(_3233_) );
	INVX1 INVX1_1092 ( .A(micro_hash_synth_2_W_25__0_), .Y(_4772_) );
	XOR2X1 XOR2X1_66 ( .A(micro_hash_synth_2_W_11__0_), .B(micro_hash_synth_2_W_16__0_), .Y(_4773_) );
	NOR2X1 NOR2X1_482 ( .A(micro_hash_synth_2_W_22__0_), .B(_4773_), .Y(_4774_) );
	OAI22X1 OAI22X1_485 ( .A(_4735__bF_buf7), .B(_4774_), .C(_4740__bF_buf4), .D(_4772_), .Y(_3244_) );
	INVX1 INVX1_1093 ( .A(micro_hash_synth_2_W_25__1_), .Y(_4775_) );
	INVX1 INVX1_1094 ( .A(micro_hash_synth_2_W_11__1_), .Y(_4776_) );
	INVX1 INVX1_1095 ( .A(micro_hash_synth_2_W_22__1_), .Y(_4777_) );
	OAI21X1 OAI21X1_1223 ( .A(_4776_), .B(micro_hash_synth_2_W_16__1_), .C(_4777_), .Y(_4778_) );
	AOI21X1 AOI21X1_854 ( .A(_4776_), .B(micro_hash_synth_2_W_16__1_), .C(_4778_), .Y(_4779_) );
	OAI22X1 OAI22X1_486 ( .A(_4735__bF_buf6), .B(_4779_), .C(_4740__bF_buf3), .D(_4775_), .Y(_3255_) );
	INVX1 INVX1_1096 ( .A(micro_hash_synth_2_W_25__2_), .Y(_4780_) );
	INVX1 INVX1_1097 ( .A(micro_hash_synth_2_W_11__2_), .Y(_4781_) );
	INVX1 INVX1_1098 ( .A(micro_hash_synth_2_W_22__2_), .Y(_4782_) );
	OAI21X1 OAI21X1_1224 ( .A(_4781_), .B(micro_hash_synth_2_W_16__2_), .C(_4782_), .Y(_4783_) );
	AOI21X1 AOI21X1_855 ( .A(_4781_), .B(micro_hash_synth_2_W_16__2_), .C(_4783_), .Y(_4784_) );
	OAI22X1 OAI22X1_487 ( .A(_4735__bF_buf5), .B(_4784_), .C(_4740__bF_buf2), .D(_4780_), .Y(_3266_) );
	INVX1 INVX1_1099 ( .A(micro_hash_synth_2_W_25__3_), .Y(_4785_) );
	XOR2X1 XOR2X1_67 ( .A(micro_hash_synth_2_W_11__3_), .B(micro_hash_synth_2_W_16__3_), .Y(_4786_) );
	NOR2X1 NOR2X1_483 ( .A(micro_hash_synth_2_W_22__3_), .B(_4786_), .Y(_4787_) );
	OAI22X1 OAI22X1_488 ( .A(_4735__bF_buf4), .B(_4787_), .C(_4740__bF_buf1), .D(_4785_), .Y(_3277_) );
	INVX1 INVX1_1100 ( .A(micro_hash_synth_2_W_25__4_), .Y(_4788_) );
	XOR2X1 XOR2X1_68 ( .A(micro_hash_synth_2_W_11__4_), .B(micro_hash_synth_2_W_16__4_), .Y(_4789_) );
	NOR2X1 NOR2X1_484 ( .A(micro_hash_synth_2_W_22__4_), .B(_4789_), .Y(_4790_) );
	OAI22X1 OAI22X1_489 ( .A(_4735__bF_buf3), .B(_4790_), .C(_4740__bF_buf0), .D(_4788_), .Y(_3288_) );
	INVX1 INVX1_1101 ( .A(micro_hash_synth_2_W_25__5_), .Y(_4791_) );
	XOR2X1 XOR2X1_69 ( .A(micro_hash_synth_2_W_11__5_), .B(micro_hash_synth_2_W_16__5_), .Y(_4792_) );
	NOR2X1 NOR2X1_485 ( .A(micro_hash_synth_2_W_22__5_), .B(_4792_), .Y(_4793_) );
	OAI22X1 OAI22X1_490 ( .A(_4735__bF_buf2), .B(_4793_), .C(_4740__bF_buf13), .D(_4791_), .Y(_3295_) );
	INVX1 INVX1_1102 ( .A(micro_hash_synth_2_W_25__6_), .Y(_4794_) );
	XOR2X1 XOR2X1_70 ( .A(micro_hash_synth_2_W_11__6_), .B(micro_hash_synth_2_W_16__6_), .Y(_4795_) );
	NOR2X1 NOR2X1_486 ( .A(micro_hash_synth_2_W_22__6_), .B(_4795_), .Y(_4796_) );
	OAI22X1 OAI22X1_491 ( .A(_4735__bF_buf1), .B(_4796_), .C(_4740__bF_buf12), .D(_4794_), .Y(_3296_) );
	INVX1 INVX1_1103 ( .A(micro_hash_synth_2_W_25__7_), .Y(_4797_) );
	XOR2X1 XOR2X1_71 ( .A(micro_hash_synth_2_W_11__7_), .B(micro_hash_synth_2_W_16__7_), .Y(_4798_) );
	NOR2X1 NOR2X1_487 ( .A(micro_hash_synth_2_W_22__7_), .B(_4798_), .Y(_4799_) );
	OAI22X1 OAI22X1_492 ( .A(_4735__bF_buf0), .B(_4799_), .C(_4740__bF_buf11), .D(_4797_), .Y(_3297_) );
	INVX1 INVX1_1104 ( .A(micro_hash_synth_2_W_8__0_), .Y(_4800_) );
	INVX1 INVX1_1105 ( .A(bloque_in_1_64_), .Y(_4801_) );
	OAI22X1 OAI22X1_493 ( .A(_4801_), .B(_4735__bF_buf15), .C(_4740__bF_buf10), .D(_4800_), .Y(_3302_) );
	INVX1 INVX1_1106 ( .A(micro_hash_synth_2_W_8__1_), .Y(_4802_) );
	INVX1 INVX1_1107 ( .A(bloque_in_1_65_), .Y(_4803_) );
	OAI22X1 OAI22X1_494 ( .A(_4803_), .B(_4735__bF_buf14), .C(_4740__bF_buf9), .D(_4802_), .Y(_3307_) );
	INVX1 INVX1_1108 ( .A(micro_hash_synth_2_W_8__2_), .Y(_4804_) );
	INVX1 INVX1_1109 ( .A(bloque_in_1_66_), .Y(_4805_) );
	OAI22X1 OAI22X1_495 ( .A(_4805_), .B(_4735__bF_buf13), .C(_4740__bF_buf8), .D(_4804_), .Y(_3308_) );
	INVX1 INVX1_1110 ( .A(micro_hash_synth_2_W_8__3_), .Y(_4806_) );
	INVX1 INVX1_1111 ( .A(bloque_in_1_67_), .Y(_4807_) );
	OAI22X1 OAI22X1_496 ( .A(_4807_), .B(_4735__bF_buf12), .C(_4740__bF_buf7), .D(_4806_), .Y(_3309_) );
	INVX1 INVX1_1112 ( .A(micro_hash_synth_2_W_8__4_), .Y(_4808_) );
	INVX1 INVX1_1113 ( .A(bloque_in_1_68_), .Y(_4809_) );
	OAI22X1 OAI22X1_497 ( .A(_4809_), .B(_4735__bF_buf11), .C(_4740__bF_buf6), .D(_4808_), .Y(_3054_) );
	INVX1 INVX1_1114 ( .A(micro_hash_synth_2_W_8__5_), .Y(_4810_) );
	INVX1 INVX1_1115 ( .A(bloque_in_1_69_), .Y(_4811_) );
	OAI22X1 OAI22X1_498 ( .A(_4811_), .B(_4735__bF_buf10), .C(_4740__bF_buf5), .D(_4810_), .Y(_3055_) );
	INVX1 INVX1_1116 ( .A(micro_hash_synth_2_W_8__6_), .Y(_4812_) );
	INVX1 INVX1_1117 ( .A(bloque_in_1_70_), .Y(_4813_) );
	OAI22X1 OAI22X1_499 ( .A(_4813_), .B(_4735__bF_buf9), .C(_4740__bF_buf4), .D(_4812_), .Y(_3063_) );
	INVX1 INVX1_1118 ( .A(micro_hash_synth_2_W_8__7_), .Y(_4814_) );
	INVX1 INVX1_1119 ( .A(bloque_in_1_71_), .Y(_4815_) );
	OAI22X1 OAI22X1_500 ( .A(_4815_), .B(_4735__bF_buf8), .C(_4740__bF_buf3), .D(_4814_), .Y(_3065_) );
	INVX1 INVX1_1120 ( .A(micro_hash_synth_2_W_3__0_), .Y(_4816_) );
	INVX1 INVX1_1121 ( .A(bloque_in_1_24_), .Y(_4817_) );
	OAI22X1 OAI22X1_501 ( .A(_4817_), .B(_4735__bF_buf7), .C(_4740__bF_buf2), .D(_4816_), .Y(_3066_) );
	INVX1 INVX1_1122 ( .A(micro_hash_synth_2_W_3__1_), .Y(_4818_) );
	INVX1 INVX1_1123 ( .A(bloque_in_1_25_), .Y(_4819_) );
	OAI22X1 OAI22X1_502 ( .A(_4819_), .B(_4735__bF_buf6), .C(_4740__bF_buf1), .D(_4818_), .Y(_3067_) );
	INVX1 INVX1_1124 ( .A(micro_hash_synth_2_W_3__2_), .Y(_4820_) );
	INVX1 INVX1_1125 ( .A(bloque_in_1_26_), .Y(_4821_) );
	OAI22X1 OAI22X1_503 ( .A(_4821_), .B(_4735__bF_buf5), .C(_4740__bF_buf0), .D(_4820_), .Y(_3076_) );
	INVX1 INVX1_1126 ( .A(micro_hash_synth_2_W_3__3_), .Y(_4822_) );
	INVX1 INVX1_1127 ( .A(bloque_in_1_27_), .Y(_4823_) );
	OAI22X1 OAI22X1_504 ( .A(_4823_), .B(_4735__bF_buf4), .C(_4740__bF_buf13), .D(_4822_), .Y(_3079_) );
	INVX1 INVX1_1128 ( .A(micro_hash_synth_2_W_3__4_), .Y(_4824_) );
	INVX1 INVX1_1129 ( .A(bloque_in_1_28_), .Y(_4825_) );
	OAI22X1 OAI22X1_505 ( .A(_4825_), .B(_4735__bF_buf3), .C(_4740__bF_buf12), .D(_4824_), .Y(_3095_) );
	INVX1 INVX1_1130 ( .A(micro_hash_synth_2_W_3__5_), .Y(_4826_) );
	INVX1 INVX1_1131 ( .A(bloque_in_1_29_), .Y(_4827_) );
	OAI22X1 OAI22X1_506 ( .A(_4827_), .B(_4735__bF_buf2), .C(_4740__bF_buf11), .D(_4826_), .Y(_3111_) );
	INVX1 INVX1_1132 ( .A(micro_hash_synth_2_W_3__6_), .Y(_4828_) );
	INVX1 INVX1_1133 ( .A(bloque_in_1_30_), .Y(_4829_) );
	OAI22X1 OAI22X1_507 ( .A(_4829_), .B(_4735__bF_buf1), .C(_4740__bF_buf10), .D(_4828_), .Y(_3127_) );
	INVX1 INVX1_1134 ( .A(micro_hash_synth_2_W_3__7_), .Y(_4830_) );
	INVX1 INVX1_1135 ( .A(bloque_in_1_31_), .Y(_4831_) );
	OAI22X1 OAI22X1_508 ( .A(_4831_), .B(_4735__bF_buf0), .C(_4740__bF_buf9), .D(_4830_), .Y(_3143_) );
	INVX8 INVX8_10 ( .A(reset_L_bF_buf48), .Y(_4832_) );
	INVX1 INVX1_1136 ( .A(micro_hash_synth_2_W_1__0_), .Y(_4833_) );
	NOR2X1 NOR2X1_488 ( .A(_4832__bF_buf4), .B(_4833_), .Y(_3052__8_) );
	INVX1 INVX1_1137 ( .A(micro_hash_synth_2_W_1__1_), .Y(_4834_) );
	NOR2X1 NOR2X1_489 ( .A(_4832__bF_buf3), .B(_4834_), .Y(_3052__9_) );
	INVX1 INVX1_1138 ( .A(micro_hash_synth_2_W_1__2_), .Y(_4835_) );
	NOR2X1 NOR2X1_490 ( .A(_4832__bF_buf2), .B(_4835_), .Y(_3052__10_) );
	INVX1 INVX1_1139 ( .A(micro_hash_synth_2_W_1__3_), .Y(_4836_) );
	NOR2X1 NOR2X1_491 ( .A(_4832__bF_buf1), .B(_4836_), .Y(_3052__11_) );
	INVX1 INVX1_1140 ( .A(micro_hash_synth_2_W_1__4_), .Y(_4837_) );
	NOR2X1 NOR2X1_492 ( .A(_4832__bF_buf0), .B(_4837_), .Y(_3052__12_) );
	INVX1 INVX1_1141 ( .A(micro_hash_synth_2_W_1__5_), .Y(_4838_) );
	NOR2X1 NOR2X1_493 ( .A(_4832__bF_buf5), .B(_4838_), .Y(_3052__13_) );
	INVX1 INVX1_1142 ( .A(micro_hash_synth_2_W_1__6_), .Y(_4839_) );
	NOR2X1 NOR2X1_494 ( .A(_4832__bF_buf4), .B(_4839_), .Y(_3052__14_) );
	INVX1 INVX1_1143 ( .A(micro_hash_synth_2_W_1__7_), .Y(_4840_) );
	NOR2X1 NOR2X1_495 ( .A(_4832__bF_buf3), .B(_4840_), .Y(_3052__15_) );
	INVX1 INVX1_1144 ( .A(micro_hash_synth_2_W_0__0_), .Y(_4841_) );
	NOR2X1 NOR2X1_496 ( .A(_4832__bF_buf2), .B(_4841_), .Y(_3052__0_) );
	INVX1 INVX1_1145 ( .A(micro_hash_synth_2_W_0__1_), .Y(_4842_) );
	NOR2X1 NOR2X1_497 ( .A(_4832__bF_buf1), .B(_4842_), .Y(_3052__1_) );
	INVX1 INVX1_1146 ( .A(micro_hash_synth_2_W_0__2_), .Y(_4843_) );
	NOR2X1 NOR2X1_498 ( .A(_4832__bF_buf0), .B(_4843_), .Y(_3052__2_) );
	INVX1 INVX1_1147 ( .A(micro_hash_synth_2_W_0__3_), .Y(_4844_) );
	NOR2X1 NOR2X1_499 ( .A(_4832__bF_buf5), .B(_4844_), .Y(_3052__3_) );
	INVX1 INVX1_1148 ( .A(micro_hash_synth_2_W_0__4_), .Y(_4845_) );
	NOR2X1 NOR2X1_500 ( .A(_4832__bF_buf4), .B(_4845_), .Y(_3052__4_) );
	INVX1 INVX1_1149 ( .A(micro_hash_synth_2_W_0__5_), .Y(_4846_) );
	NOR2X1 NOR2X1_501 ( .A(_4832__bF_buf3), .B(_4846_), .Y(_3052__5_) );
	INVX1 INVX1_1150 ( .A(micro_hash_synth_2_W_0__6_), .Y(_4847_) );
	NOR2X1 NOR2X1_502 ( .A(_4832__bF_buf2), .B(_4847_), .Y(_3052__6_) );
	INVX1 INVX1_1151 ( .A(micro_hash_synth_2_W_0__7_), .Y(_4848_) );
	NOR2X1 NOR2X1_503 ( .A(_4832__bF_buf1), .B(_4848_), .Y(_3052__7_) );
	INVX1 INVX1_1152 ( .A(micro_hash_synth_2_W_2__0_), .Y(_4849_) );
	NOR2X1 NOR2X1_504 ( .A(_4832__bF_buf0), .B(_4849_), .Y(_3052__16_) );
	INVX1 INVX1_1153 ( .A(micro_hash_synth_2_W_2__1_), .Y(_4850_) );
	NOR2X1 NOR2X1_505 ( .A(_4832__bF_buf5), .B(_4850_), .Y(_3052__17_) );
	INVX1 INVX1_1154 ( .A(micro_hash_synth_2_W_2__2_), .Y(_4851_) );
	NOR2X1 NOR2X1_506 ( .A(_4832__bF_buf4), .B(_4851_), .Y(_3052__18_) );
	INVX1 INVX1_1155 ( .A(micro_hash_synth_2_W_2__3_), .Y(_4852_) );
	NOR2X1 NOR2X1_507 ( .A(_4832__bF_buf3), .B(_4852_), .Y(_3052__19_) );
	INVX1 INVX1_1156 ( .A(micro_hash_synth_2_W_2__4_), .Y(_4853_) );
	NOR2X1 NOR2X1_508 ( .A(_4832__bF_buf2), .B(_4853_), .Y(_3052__20_) );
	INVX1 INVX1_1157 ( .A(micro_hash_synth_2_W_2__5_), .Y(_4854_) );
	NOR2X1 NOR2X1_509 ( .A(_4832__bF_buf1), .B(_4854_), .Y(_3052__21_) );
	INVX1 INVX1_1158 ( .A(micro_hash_synth_2_W_2__6_), .Y(_4855_) );
	NOR2X1 NOR2X1_510 ( .A(_4832__bF_buf0), .B(_4855_), .Y(_3052__22_) );
	INVX1 INVX1_1159 ( .A(micro_hash_synth_2_W_2__7_), .Y(_4856_) );
	NOR2X1 NOR2X1_511 ( .A(_4832__bF_buf5), .B(_4856_), .Y(_3052__23_) );
	NOR2X1 NOR2X1_512 ( .A(_4832__bF_buf4), .B(_4816_), .Y(_3052__24_) );
	NOR2X1 NOR2X1_513 ( .A(_4832__bF_buf3), .B(_4818_), .Y(_3052__25_) );
	NOR2X1 NOR2X1_514 ( .A(_4832__bF_buf2), .B(_4820_), .Y(_3052__26_) );
	NOR2X1 NOR2X1_515 ( .A(_4832__bF_buf1), .B(_4822_), .Y(_3052__27_) );
	NOR2X1 NOR2X1_516 ( .A(_4832__bF_buf0), .B(_4824_), .Y(_3052__28_) );
	NOR2X1 NOR2X1_517 ( .A(_4832__bF_buf5), .B(_4826_), .Y(_3052__29_) );
	NOR2X1 NOR2X1_518 ( .A(_4832__bF_buf4), .B(_4828_), .Y(_3052__30_) );
	NOR2X1 NOR2X1_519 ( .A(_4832__bF_buf3), .B(_4830_), .Y(_3052__31_) );
	INVX1 INVX1_1160 ( .A(Hhash_synth2_8_), .Y(_3310_) );
	NOR2X1 NOR2X1_520 ( .A(concatenador_counter_2d_4_), .B(_4737_), .Y(_3311_) );
	INVX1 INVX1_1161 ( .A(_3311_), .Y(_3312_) );
	INVX1 INVX1_1162 ( .A(concatenador_counter_2d_5_), .Y(_3313_) );
	NOR2X1 NOR2X1_521 ( .A(_1__bF_buf1), .B(_3313_), .Y(_3314_) );
	NAND2X1 NAND2X1_661 ( .A(concatenador_counter_2d_0_bF_buf6), .B(_3314_), .Y(_3315_) );
	NOR2X1 NOR2X1_522 ( .A(_3315_), .B(_3312_), .Y(_3316_) );
	INVX2 INVX2_9 ( .A(_3316__bF_buf2), .Y(_3317_) );
	NOR2X1 NOR2X1_523 ( .A(_4832__bF_buf2), .B(_3317_), .Y(_3318_) );
	NAND3X1 NAND3X1_216 ( .A(reset_L_bF_buf47), .B(_4739_), .C(_3317_), .Y(_3319_) );
	INVX4 INVX4_8 ( .A(_3318_), .Y(_3320_) );
	OAI21X1 OAI21X1_1225 ( .A(_3320_), .B(micro_hash_synth_2_b_0_), .C(_3319_), .Y(_3321_) );
	INVX1 INVX1_1163 ( .A(micro_hash_synth_2_b_0_), .Y(_3322_) );
	NOR2X1 NOR2X1_524 ( .A(_3310_), .B(_3322_), .Y(_3323_) );
	AOI22X1 AOI22X1_37 ( .A(_3318_), .B(_3323_), .C(_3321_), .D(_3310_), .Y(_3047__8_) );
	INVX1 INVX1_1164 ( .A(Hhash_synth2_9_), .Y(_3324_) );
	INVX1 INVX1_1165 ( .A(micro_hash_synth_2_b_1_), .Y(_3325_) );
	NOR2X1 NOR2X1_525 ( .A(_3324_), .B(_3325_), .Y(_3326_) );
	NOR2X1 NOR2X1_526 ( .A(Hhash_synth2_9_), .B(micro_hash_synth_2_b_1_), .Y(_3327_) );
	NOR2X1 NOR2X1_527 ( .A(_3327_), .B(_3326_), .Y(_3328_) );
	NAND2X1 NAND2X1_662 ( .A(_3323_), .B(_3328_), .Y(_3329_) );
	OR2X2 OR2X2_58 ( .A(_3328_), .B(_3323_), .Y(_3330_) );
	AOI21X1 AOI21X1_856 ( .A(_3329_), .B(_3330_), .C(_3317_), .Y(_3331_) );
	OAI21X1 OAI21X1_1226 ( .A(_4737_), .B(_4731_), .C(reset_L_bF_buf46), .Y(_3332_) );
	INVX4 INVX4_9 ( .A(_3332__bF_buf3), .Y(_3333_) );
	NAND2X1 NAND2X1_663 ( .A(Hhash_synth2_9_), .B(_3333__bF_buf3), .Y(_3334_) );
	AOI21X1 AOI21X1_857 ( .A(_3334_), .B(_3320_), .C(_3331_), .Y(_3047__9_) );
	OAI21X1 OAI21X1_1227 ( .A(_3324_), .B(_3325_), .C(_3329_), .Y(_3335_) );
	AND2X2 AND2X2_92 ( .A(Hhash_synth2_10_), .B(micro_hash_synth_2_b_2_), .Y(_3336_) );
	NOR2X1 NOR2X1_528 ( .A(Hhash_synth2_10_), .B(micro_hash_synth_2_b_2_), .Y(_3337_) );
	NOR2X1 NOR2X1_529 ( .A(_3337_), .B(_3336_), .Y(_3338_) );
	XNOR2X1 XNOR2X1_48 ( .A(_3335_), .B(_3338_), .Y(_3339_) );
	NAND2X1 NAND2X1_664 ( .A(Hhash_synth2_10_), .B(_3333__bF_buf2), .Y(_3340_) );
	AOI22X1 AOI22X1_38 ( .A(_3316__bF_buf1), .B(_3339_), .C(_3320_), .D(_3340_), .Y(_3047__10_) );
	AOI21X1 AOI21X1_858 ( .A(_3338_), .B(_3335_), .C(_3336_), .Y(_3341_) );
	INVX1 INVX1_1166 ( .A(Hhash_synth2_11_), .Y(_3342_) );
	INVX1 INVX1_1167 ( .A(micro_hash_synth_2_b_3_), .Y(_3343_) );
	NOR2X1 NOR2X1_530 ( .A(_3342_), .B(_3343_), .Y(_3344_) );
	NOR2X1 NOR2X1_531 ( .A(Hhash_synth2_11_), .B(micro_hash_synth_2_b_3_), .Y(_3345_) );
	NOR2X1 NOR2X1_532 ( .A(_3345_), .B(_3344_), .Y(_3346_) );
	XOR2X1 XOR2X1_72 ( .A(_3341_), .B(_3346_), .Y(_3347_) );
	OAI21X1 OAI21X1_1228 ( .A(Hhash_synth2_11_), .B(_3332__bF_buf2), .C(_3320_), .Y(_3348_) );
	OAI21X1 OAI21X1_1229 ( .A(_3317_), .B(_3347_), .C(_3348_), .Y(_3047__11_) );
	XOR2X1 XOR2X1_73 ( .A(Hhash_synth2_12_), .B(micro_hash_synth_2_b_4_), .Y(_3349_) );
	INVX1 INVX1_1168 ( .A(_3344_), .Y(_3350_) );
	OAI21X1 OAI21X1_1230 ( .A(_3341_), .B(_3345_), .C(_3350_), .Y(_3351_) );
	XNOR2X1 XNOR2X1_49 ( .A(_3351_), .B(_3349_), .Y(_3352_) );
	AOI21X1 AOI21X1_859 ( .A(Hhash_synth2_12_), .B(_3333__bF_buf1), .C(_3318_), .Y(_3353_) );
	AOI21X1 AOI21X1_860 ( .A(_3316__bF_buf0), .B(_3352_), .C(_3353_), .Y(_3047__12_) );
	AOI21X1 AOI21X1_861 ( .A(Hhash_synth2_13_), .B(_3333__bF_buf0), .C(_3318_), .Y(_3354_) );
	AND2X2 AND2X2_93 ( .A(_3351_), .B(_3349_), .Y(_3355_) );
	AOI21X1 AOI21X1_862 ( .A(Hhash_synth2_12_), .B(micro_hash_synth_2_b_4_), .C(_3355_), .Y(_3356_) );
	NAND2X1 NAND2X1_665 ( .A(Hhash_synth2_13_), .B(micro_hash_synth_2_b_5_), .Y(_3357_) );
	INVX1 INVX1_1169 ( .A(_3357_), .Y(_3358_) );
	NOR2X1 NOR2X1_533 ( .A(Hhash_synth2_13_), .B(micro_hash_synth_2_b_5_), .Y(_3359_) );
	NOR2X1 NOR2X1_534 ( .A(_3359_), .B(_3358_), .Y(_3360_) );
	XOR2X1 XOR2X1_74 ( .A(_3356_), .B(_3360_), .Y(_3361_) );
	AOI21X1 AOI21X1_863 ( .A(_3316__bF_buf3), .B(_3361_), .C(_3354_), .Y(_3047__13_) );
	XOR2X1 XOR2X1_75 ( .A(Hhash_synth2_14_), .B(micro_hash_synth_2_b_6_), .Y(_3362_) );
	OAI21X1 OAI21X1_1231 ( .A(_3356_), .B(_3359_), .C(_3357_), .Y(_3363_) );
	XNOR2X1 XNOR2X1_50 ( .A(_3363_), .B(_3362_), .Y(_3364_) );
	AOI21X1 AOI21X1_864 ( .A(Hhash_synth2_14_), .B(_3333__bF_buf3), .C(_3318_), .Y(_3365_) );
	AOI21X1 AOI21X1_865 ( .A(_3316__bF_buf2), .B(_3364_), .C(_3365_), .Y(_3047__14_) );
	OAI21X1 OAI21X1_1232 ( .A(Hhash_synth2_15_), .B(_3332__bF_buf1), .C(_3320_), .Y(_3366_) );
	AND2X2 AND2X2_94 ( .A(Hhash_synth2_14_), .B(micro_hash_synth_2_b_6_), .Y(_3367_) );
	AOI21X1 AOI21X1_866 ( .A(_3362_), .B(_3363_), .C(_3367_), .Y(_3368_) );
	XNOR2X1 XNOR2X1_51 ( .A(Hhash_synth2_15_), .B(micro_hash_synth_2_b_7_), .Y(_3369_) );
	NOR2X1 NOR2X1_535 ( .A(_3369_), .B(_3368_), .Y(_3370_) );
	NAND2X1 NAND2X1_666 ( .A(_3369_), .B(_3368_), .Y(_3371_) );
	NAND2X1 NAND2X1_667 ( .A(_3316__bF_buf1), .B(_3371_), .Y(_3372_) );
	OAI21X1 OAI21X1_1233 ( .A(_3372_), .B(_3370_), .C(_3366_), .Y(_3047__15_) );
	INVX1 INVX1_1170 ( .A(Hhash_synth2_0_), .Y(_3373_) );
	OAI21X1 OAI21X1_1234 ( .A(_3320_), .B(micro_hash_synth_2_a_0_), .C(_3319_), .Y(_3374_) );
	INVX1 INVX1_1171 ( .A(micro_hash_synth_2_a_0_), .Y(_3375_) );
	NOR2X1 NOR2X1_536 ( .A(_3373_), .B(_3375_), .Y(_3376_) );
	AOI22X1 AOI22X1_39 ( .A(_3318_), .B(_3376_), .C(_3374_), .D(_3373_), .Y(_3047__0_) );
	INVX1 INVX1_1172 ( .A(Hhash_synth2_1_), .Y(_3377_) );
	INVX1 INVX1_1173 ( .A(micro_hash_synth_2_a_1_), .Y(_3378_) );
	NOR2X1 NOR2X1_537 ( .A(_3377_), .B(_3378_), .Y(_3379_) );
	NOR2X1 NOR2X1_538 ( .A(Hhash_synth2_1_), .B(micro_hash_synth_2_a_1_), .Y(_3380_) );
	NOR2X1 NOR2X1_539 ( .A(_3380_), .B(_3379_), .Y(_3381_) );
	NAND2X1 NAND2X1_668 ( .A(_3376_), .B(_3381_), .Y(_3382_) );
	OR2X2 OR2X2_59 ( .A(_3381_), .B(_3376_), .Y(_3383_) );
	AOI21X1 AOI21X1_867 ( .A(_3382_), .B(_3383_), .C(_3317_), .Y(_3384_) );
	NAND2X1 NAND2X1_669 ( .A(Hhash_synth2_1_), .B(_3333__bF_buf2), .Y(_3385_) );
	AOI21X1 AOI21X1_868 ( .A(_3385_), .B(_3320_), .C(_3384_), .Y(_3047__1_) );
	OAI21X1 OAI21X1_1235 ( .A(_3377_), .B(_3378_), .C(_3382_), .Y(_3386_) );
	AND2X2 AND2X2_95 ( .A(Hhash_synth2_2_), .B(micro_hash_synth_2_a_2_), .Y(_3387_) );
	NOR2X1 NOR2X1_540 ( .A(Hhash_synth2_2_), .B(micro_hash_synth_2_a_2_), .Y(_3388_) );
	NOR2X1 NOR2X1_541 ( .A(_3388_), .B(_3387_), .Y(_3389_) );
	XNOR2X1 XNOR2X1_52 ( .A(_3386_), .B(_3389_), .Y(_3390_) );
	NAND2X1 NAND2X1_670 ( .A(Hhash_synth2_2_), .B(_3333__bF_buf1), .Y(_3391_) );
	AOI22X1 AOI22X1_40 ( .A(_3316__bF_buf0), .B(_3390_), .C(_3320_), .D(_3391_), .Y(_3047__2_) );
	NAND2X1 NAND2X1_671 ( .A(Hhash_synth2_3_), .B(_3333__bF_buf0), .Y(_3392_) );
	AOI21X1 AOI21X1_869 ( .A(_3389_), .B(_3386_), .C(_3387_), .Y(_3393_) );
	AND2X2 AND2X2_96 ( .A(Hhash_synth2_3_), .B(micro_hash_synth_2_a_3_), .Y(_3394_) );
	NOR2X1 NOR2X1_542 ( .A(Hhash_synth2_3_), .B(micro_hash_synth_2_a_3_), .Y(_3395_) );
	NOR2X1 NOR2X1_543 ( .A(_3395_), .B(_3394_), .Y(_3396_) );
	XOR2X1 XOR2X1_76 ( .A(_3393_), .B(_3396_), .Y(_3397_) );
	AOI22X1 AOI22X1_41 ( .A(_3316__bF_buf3), .B(_3397_), .C(_3320_), .D(_3392_), .Y(_3047__3_) );
	XOR2X1 XOR2X1_77 ( .A(Hhash_synth2_4_), .B(micro_hash_synth_2_a_4_), .Y(_3398_) );
	INVX1 INVX1_1174 ( .A(_3394_), .Y(_3399_) );
	OAI21X1 OAI21X1_1236 ( .A(_3393_), .B(_3395_), .C(_3399_), .Y(_3400_) );
	XNOR2X1 XNOR2X1_53 ( .A(_3400_), .B(_3398_), .Y(_3401_) );
	AOI21X1 AOI21X1_870 ( .A(Hhash_synth2_4_), .B(_3333__bF_buf3), .C(_3318_), .Y(_3402_) );
	AOI21X1 AOI21X1_871 ( .A(_3316__bF_buf2), .B(_3401_), .C(_3402_), .Y(_3047__4_) );
	AOI21X1 AOI21X1_872 ( .A(Hhash_synth2_5_), .B(_3333__bF_buf2), .C(_3318_), .Y(_3403_) );
	AND2X2 AND2X2_97 ( .A(_3400_), .B(_3398_), .Y(_3404_) );
	AOI21X1 AOI21X1_873 ( .A(Hhash_synth2_4_), .B(micro_hash_synth_2_a_4_), .C(_3404_), .Y(_3405_) );
	NAND2X1 NAND2X1_672 ( .A(Hhash_synth2_5_), .B(micro_hash_synth_2_a_5_), .Y(_3406_) );
	INVX1 INVX1_1175 ( .A(_3406_), .Y(_3407_) );
	NOR2X1 NOR2X1_544 ( .A(Hhash_synth2_5_), .B(micro_hash_synth_2_a_5_), .Y(_3408_) );
	NOR2X1 NOR2X1_545 ( .A(_3408_), .B(_3407_), .Y(_3409_) );
	OAI21X1 OAI21X1_1237 ( .A(_3405_), .B(_3409_), .C(_3316__bF_buf1), .Y(_3410_) );
	AOI21X1 AOI21X1_874 ( .A(_3405_), .B(_3409_), .C(_3410_), .Y(_3411_) );
	NOR2X1 NOR2X1_546 ( .A(_3403_), .B(_3411_), .Y(_3047__5_) );
	XOR2X1 XOR2X1_78 ( .A(Hhash_synth2_6_), .B(micro_hash_synth_2_a_6_), .Y(_3412_) );
	OAI21X1 OAI21X1_1238 ( .A(_3405_), .B(_3408_), .C(_3406_), .Y(_3413_) );
	XNOR2X1 XNOR2X1_54 ( .A(_3413_), .B(_3412_), .Y(_3414_) );
	AOI21X1 AOI21X1_875 ( .A(Hhash_synth2_6_), .B(_3333__bF_buf1), .C(_3318_), .Y(_3415_) );
	AOI21X1 AOI21X1_876 ( .A(_3316__bF_buf0), .B(_3414_), .C(_3415_), .Y(_3047__6_) );
	AOI21X1 AOI21X1_877 ( .A(Hhash_synth2_7_), .B(_3333__bF_buf0), .C(_3318_), .Y(_3416_) );
	INVX1 INVX1_1176 ( .A(Hhash_synth2_6_), .Y(_3417_) );
	INVX1 INVX1_1177 ( .A(micro_hash_synth_2_a_6_), .Y(_3418_) );
	NAND2X1 NAND2X1_673 ( .A(_3412_), .B(_3413_), .Y(_3419_) );
	OAI21X1 OAI21X1_1239 ( .A(_3417_), .B(_3418_), .C(_3419_), .Y(_3420_) );
	XNOR2X1 XNOR2X1_55 ( .A(Hhash_synth2_7_), .B(micro_hash_synth_2_a_7_), .Y(_3421_) );
	OAI21X1 OAI21X1_1240 ( .A(_3420_), .B(_3421_), .C(_3316__bF_buf3), .Y(_3422_) );
	AOI21X1 AOI21X1_878 ( .A(_3420_), .B(_3421_), .C(_3422_), .Y(_3423_) );
	NOR2X1 NOR2X1_547 ( .A(_3416_), .B(_3423_), .Y(_3047__7_) );
	OAI21X1 OAI21X1_1241 ( .A(_4737_), .B(concatenador_counter_2d_4_), .C(concatenador_counter_2d_5_), .Y(_3424_) );
	NOR2X1 NOR2X1_548 ( .A(_4832__bF_buf1), .B(_3424__bF_buf1), .Y(_3425_) );
	INVX4 INVX4_10 ( .A(_3425_), .Y(_3426_) );
	OR2X2 OR2X2_60 ( .A(_3426_), .B(micro_hash_synth_2_k_0_), .Y(_3051__0_) );
	INVX1 INVX1_1178 ( .A(micro_hash_synth_2_k_1_), .Y(_3427_) );
	NOR2X1 NOR2X1_549 ( .A(_3427_), .B(_3426_), .Y(_3051__1_) );
	INVX1 INVX1_1179 ( .A(micro_hash_synth_2_k_2_), .Y(_3428_) );
	NOR2X1 NOR2X1_550 ( .A(_3428_), .B(_3426_), .Y(_3051__2_) );
	INVX1 INVX1_1180 ( .A(micro_hash_synth_2_k_3_), .Y(_3429_) );
	NOR2X1 NOR2X1_551 ( .A(concatenador_counter_2d_0_bF_buf5), .B(concatenador_counter_2d_5_), .Y(_3430_) );
	AOI21X1 AOI21X1_879 ( .A(_3430_), .B(_4736_), .C(_4730_), .Y(_3431_) );
	INVX1 INVX1_1181 ( .A(_3431_), .Y(_3432_) );
	NOR2X1 NOR2X1_552 ( .A(_4832__bF_buf0), .B(_3432_), .Y(_3433_) );
	OAI21X1 OAI21X1_1242 ( .A(_3424__bF_buf0), .B(_3429_), .C(_3433_), .Y(_3051__3_) );
	INVX1 INVX1_1182 ( .A(micro_hash_synth_2_k_4_), .Y(_3434_) );
	OAI21X1 OAI21X1_1243 ( .A(_3424__bF_buf3), .B(_3434_), .C(_3433_), .Y(_3051__4_) );
	INVX1 INVX1_1183 ( .A(micro_hash_synth_2_k_5_), .Y(_3435_) );
	INVX2 INVX2_10 ( .A(_3424__bF_buf2), .Y(_3436_) );
	INVX2 INVX2_11 ( .A(_3433_), .Y(_3437_) );
	AOI21X1 AOI21X1_880 ( .A(_3435_), .B(_3436_), .C(_3437_), .Y(_3051__5_) );
	AND2X2 AND2X2_98 ( .A(_3425_), .B(micro_hash_synth_2_k_6_), .Y(_3051__6_) );
	OR2X2 OR2X2_61 ( .A(_3426_), .B(micro_hash_synth_2_k_7_), .Y(_3051__7_) );
	INVX1 INVX1_1184 ( .A(micro_hash_synth_2_c_0_), .Y(_3438_) );
	INVX4 INVX4_11 ( .A(concatenador_counter_2d_1_bF_buf4), .Y(_3439_) );
	NOR2X1 NOR2X1_553 ( .A(concatenador_counter_2d_2_), .B(_3439__bF_buf1), .Y(_3440_) );
	INVX1 INVX1_1185 ( .A(concatenador_counter_2d_2_), .Y(_3441_) );
	NOR2X1 NOR2X1_554 ( .A(concatenador_counter_2d_1_bF_buf3), .B(_3441_), .Y(_3442_) );
	NOR2X1 NOR2X1_555 ( .A(_3440__bF_buf4), .B(_3442__bF_buf2), .Y(_3443_) );
	NOR2X1 NOR2X1_556 ( .A(micro_hash_synth_2_W_5__0_), .B(_4733__bF_buf1), .Y(_3444_) );
	OAI21X1 OAI21X1_1244 ( .A(concatenador_counter_2d_0_bF_buf4), .B(micro_hash_synth_2_W_4__0_), .C(concatenador_counter_2d_1_bF_buf2), .Y(_3445_) );
	NOR2X1 NOR2X1_557 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_6__0_), .Y(_3446_) );
	OAI21X1 OAI21X1_1245 ( .A(_4733__bF_buf0), .B(micro_hash_synth_2_W_7__0_), .C(_3439__bF_buf0), .Y(_3447_) );
	OAI22X1 OAI22X1_509 ( .A(_3444_), .B(_3445_), .C(_3447_), .D(_3446_), .Y(_3448_) );
	NAND2X1 NAND2X1_674 ( .A(_3443__bF_buf5), .B(_3448_), .Y(_3449_) );
	NAND3X1 NAND3X1_217 ( .A(concatenador_counter_2d_3_), .B(_3439__bF_buf3), .C(_3441_), .Y(_3450_) );
	INVX1 INVX1_1186 ( .A(concatenador_counter_2d_3_), .Y(_3451_) );
	OAI21X1 OAI21X1_1246 ( .A(concatenador_counter_2d_1_bF_buf1), .B(concatenador_counter_2d_2_), .C(_3451_), .Y(_3452_) );
	NAND2X1 NAND2X1_675 ( .A(_3452_), .B(_3450_), .Y(_3453_) );
	NAND2X1 NAND2X1_676 ( .A(concatenador_counter_2d_0_bF_buf2), .B(micro_hash_synth_2_W_1__0_), .Y(_3454_) );
	OAI21X1 OAI21X1_1247 ( .A(_4841_), .B(concatenador_counter_2d_0_bF_buf1), .C(_3454_), .Y(_3455_) );
	NAND2X1 NAND2X1_677 ( .A(concatenador_counter_2d_0_bF_buf0), .B(micro_hash_synth_2_W_3__0_), .Y(_3456_) );
	OAI21X1 OAI21X1_1248 ( .A(_4849_), .B(concatenador_counter_2d_0_bF_buf12), .C(_3456_), .Y(_3457_) );
	AOI22X1 AOI22X1_42 ( .A(_3455_), .B(_3440__bF_buf3), .C(_3442__bF_buf1), .D(_3457_), .Y(_3458_) );
	NAND3X1 NAND3X1_218 ( .A(_3453__bF_buf0), .B(_3458_), .C(_3449_), .Y(_3459_) );
	XOR2X1 XOR2X1_79 ( .A(_4736_), .B(concatenador_counter_2d_4_), .Y(_3460_) );
	NOR2X1 NOR2X1_558 ( .A(micro_hash_synth_2_W_13__0_), .B(_4733__bF_buf7), .Y(_3461_) );
	OAI21X1 OAI21X1_1249 ( .A(concatenador_counter_2d_0_bF_buf11), .B(micro_hash_synth_2_W_12__0_), .C(concatenador_counter_2d_1_bF_buf0), .Y(_3462_) );
	NOR2X1 NOR2X1_559 ( .A(concatenador_counter_2d_0_bF_buf10), .B(micro_hash_synth_2_W_14__0_), .Y(_3463_) );
	OAI21X1 OAI21X1_1250 ( .A(_4733__bF_buf6), .B(micro_hash_synth_2_W_15__0_), .C(_3439__bF_buf2), .Y(_3464_) );
	OAI22X1 OAI22X1_510 ( .A(_3461_), .B(_3462_), .C(_3464_), .D(_3463_), .Y(_3465_) );
	NAND2X1 NAND2X1_678 ( .A(_3443__bF_buf4), .B(_3465_), .Y(_3466_) );
	NAND2X1 NAND2X1_679 ( .A(concatenador_counter_2d_1_bF_buf6), .B(_3441_), .Y(_3467_) );
	NAND2X1 NAND2X1_680 ( .A(concatenador_counter_2d_2_), .B(_3439__bF_buf1), .Y(_3468_) );
	MUX2X1 MUX2X1_39 ( .A(micro_hash_synth_2_W_11__0_), .B(micro_hash_synth_2_W_10__0_), .S(concatenador_counter_2d_0_bF_buf9), .Y(_3469_) );
	MUX2X1 MUX2X1_40 ( .A(micro_hash_synth_2_W_9__0_), .B(micro_hash_synth_2_W_8__0_), .S(concatenador_counter_2d_0_bF_buf8), .Y(_3470_) );
	OAI22X1 OAI22X1_511 ( .A(_3469_), .B(_3468_), .C(_3467_), .D(_3470_), .Y(_3471_) );
	NOR2X1 NOR2X1_560 ( .A(_3453__bF_buf3), .B(_3471_), .Y(_3472_) );
	AOI21X1 AOI21X1_881 ( .A(_3466_), .B(_3472_), .C(_3460_), .Y(_3473_) );
	NOR2X1 NOR2X1_561 ( .A(micro_hash_synth_2_W_21__0_), .B(_4733__bF_buf5), .Y(_3474_) );
	OAI21X1 OAI21X1_1251 ( .A(concatenador_counter_2d_0_bF_buf7), .B(micro_hash_synth_2_W_20__0_), .C(concatenador_counter_2d_1_bF_buf5), .Y(_3475_) );
	NOR2X1 NOR2X1_562 ( .A(concatenador_counter_2d_0_bF_buf6), .B(micro_hash_synth_2_W_22__0_), .Y(_3476_) );
	OAI21X1 OAI21X1_1252 ( .A(_4733__bF_buf4), .B(micro_hash_synth_2_W_23__0_), .C(_3439__bF_buf0), .Y(_3477_) );
	OAI22X1 OAI22X1_512 ( .A(_3474_), .B(_3475_), .C(_3477_), .D(_3476_), .Y(_3478_) );
	NAND2X1 NAND2X1_681 ( .A(_3443__bF_buf3), .B(_3478_), .Y(_3479_) );
	INVX1 INVX1_1187 ( .A(micro_hash_synth_2_W_18__0_), .Y(_3480_) );
	NAND2X1 NAND2X1_682 ( .A(concatenador_counter_2d_0_bF_buf5), .B(micro_hash_synth_2_W_19__0_), .Y(_3481_) );
	OAI21X1 OAI21X1_1253 ( .A(_3480_), .B(concatenador_counter_2d_0_bF_buf4), .C(_3481_), .Y(_3482_) );
	INVX1 INVX1_1188 ( .A(micro_hash_synth_2_W_16__0_), .Y(_3483_) );
	NAND2X1 NAND2X1_683 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_17__0_), .Y(_3484_) );
	OAI21X1 OAI21X1_1254 ( .A(_3483_), .B(concatenador_counter_2d_0_bF_buf2), .C(_3484_), .Y(_3485_) );
	AOI22X1 AOI22X1_43 ( .A(_3482_), .B(_3442__bF_buf0), .C(_3440__bF_buf2), .D(_3485_), .Y(_3486_) );
	NAND3X1 NAND3X1_219 ( .A(_3453__bF_buf2), .B(_3486_), .C(_3479_), .Y(_3487_) );
	OAI21X1 OAI21X1_1255 ( .A(concatenador_counter_2d_1_bF_buf4), .B(concatenador_counter_2d_2_), .C(concatenador_counter_2d_3_), .Y(_3488_) );
	OAI21X1 OAI21X1_1256 ( .A(_4729_), .B(concatenador_counter_2d_1_bF_buf3), .C(_3488_), .Y(_3489_) );
	XNOR2X1 XNOR2X1_56 ( .A(_4736_), .B(concatenador_counter_2d_4_), .Y(_3490_) );
	MUX2X1 MUX2X1_41 ( .A(micro_hash_synth_2_W_29__0_), .B(micro_hash_synth_2_W_28__0_), .S(concatenador_counter_2d_0_bF_buf1), .Y(_3491_) );
	MUX2X1 MUX2X1_42 ( .A(micro_hash_synth_2_W_31__0_), .B(micro_hash_synth_2_W_30__0_), .S(concatenador_counter_2d_0_bF_buf0), .Y(_3492_) );
	MUX2X1 MUX2X1_43 ( .A(_3492_), .B(_3491_), .S(_3439__bF_buf3), .Y(_3493_) );
	MUX2X1 MUX2X1_44 ( .A(micro_hash_synth_2_W_25__0_), .B(micro_hash_synth_2_W_24__0_), .S(concatenador_counter_2d_0_bF_buf12), .Y(_3494_) );
	MUX2X1 MUX2X1_45 ( .A(micro_hash_synth_2_W_27__0_), .B(micro_hash_synth_2_W_26__0_), .S(concatenador_counter_2d_0_bF_buf11), .Y(_3495_) );
	OAI22X1 OAI22X1_513 ( .A(_3494_), .B(_3467_), .C(_3468_), .D(_3495_), .Y(_3496_) );
	AOI21X1 AOI21X1_882 ( .A(_3443__bF_buf2), .B(_3493_), .C(_3496_), .Y(_3497_) );
	AOI21X1 AOI21X1_883 ( .A(_3489__bF_buf0), .B(_3497_), .C(_3490_), .Y(_3498_) );
	AOI22X1 AOI22X1_44 ( .A(_3473_), .B(_3459_), .C(_3498_), .D(_3487_), .Y(_3499_) );
	INVX1 INVX1_1189 ( .A(_3499_), .Y(_3500_) );
	NAND2X1 NAND2X1_684 ( .A(micro_hash_synth_2_k_0_), .B(micro_hash_synth_2_x_0_), .Y(_3501_) );
	INVX1 INVX1_1190 ( .A(_3501_), .Y(_3502_) );
	NOR2X1 NOR2X1_563 ( .A(micro_hash_synth_2_k_0_), .B(micro_hash_synth_2_x_0_), .Y(_3503_) );
	NOR2X1 NOR2X1_564 ( .A(_3503_), .B(_3502_), .Y(_3504_) );
	OAI21X1 OAI21X1_1257 ( .A(_4737_), .B(_4731_), .C(_3424__bF_buf1), .Y(_3505_) );
	AOI21X1 AOI21X1_884 ( .A(_3504_), .B(_3500_), .C(_3505_), .Y(_3506_) );
	OAI21X1 OAI21X1_1258 ( .A(_3500_), .B(_3504_), .C(_3506_), .Y(_3507_) );
	OAI22X1 OAI22X1_514 ( .A(_3438_), .B(_3426_), .C(_3507_), .D(_4832__bF_buf5), .Y(_3050__0_) );
	OAI21X1 OAI21X1_1259 ( .A(_3499_), .B(_3503_), .C(_3501_), .Y(_3508_) );
	NOR2X1 NOR2X1_565 ( .A(micro_hash_synth_2_W_21__1_), .B(_4733__bF_buf3), .Y(_3509_) );
	OAI21X1 OAI21X1_1260 ( .A(concatenador_counter_2d_0_bF_buf10), .B(micro_hash_synth_2_W_20__1_), .C(concatenador_counter_2d_1_bF_buf2), .Y(_3510_) );
	MUX2X1 MUX2X1_46 ( .A(micro_hash_synth_2_W_23__1_), .B(micro_hash_synth_2_W_22__1_), .S(concatenador_counter_2d_0_bF_buf9), .Y(_3511_) );
	OAI22X1 OAI22X1_515 ( .A(_3511_), .B(concatenador_counter_2d_1_bF_buf1), .C(_3509_), .D(_3510_), .Y(_3512_) );
	INVX1 INVX1_1191 ( .A(micro_hash_synth_2_W_18__1_), .Y(_3513_) );
	NAND2X1 NAND2X1_685 ( .A(concatenador_counter_2d_0_bF_buf8), .B(micro_hash_synth_2_W_19__1_), .Y(_3514_) );
	OAI21X1 OAI21X1_1261 ( .A(_3513_), .B(concatenador_counter_2d_0_bF_buf7), .C(_3514_), .Y(_3515_) );
	NAND2X1 NAND2X1_686 ( .A(_3442__bF_buf4), .B(_3515_), .Y(_3516_) );
	INVX1 INVX1_1192 ( .A(micro_hash_synth_2_W_16__1_), .Y(_3517_) );
	NAND2X1 NAND2X1_687 ( .A(concatenador_counter_2d_0_bF_buf6), .B(micro_hash_synth_2_W_17__1_), .Y(_3518_) );
	OAI21X1 OAI21X1_1262 ( .A(_3517_), .B(concatenador_counter_2d_0_bF_buf5), .C(_3518_), .Y(_3519_) );
	NAND2X1 NAND2X1_688 ( .A(_3440__bF_buf1), .B(_3519_), .Y(_3520_) );
	NAND3X1 NAND3X1_220 ( .A(_3453__bF_buf1), .B(_3516_), .C(_3520_), .Y(_3521_) );
	AOI21X1 AOI21X1_885 ( .A(_3443__bF_buf1), .B(_3512_), .C(_3521_), .Y(_3522_) );
	NAND2X1 NAND2X1_689 ( .A(_3467_), .B(_3468_), .Y(_3523_) );
	INVX1 INVX1_1193 ( .A(micro_hash_synth_2_W_29__1_), .Y(_3524_) );
	NAND2X1 NAND2X1_690 ( .A(concatenador_counter_2d_0_bF_buf4), .B(_3524_), .Y(_3525_) );
	OR2X2 OR2X2_62 ( .A(concatenador_counter_2d_0_bF_buf3), .B(micro_hash_synth_2_W_28__1_), .Y(_3526_) );
	NAND3X1 NAND3X1_221 ( .A(concatenador_counter_2d_1_bF_buf0), .B(_3526_), .C(_3525_), .Y(_3527_) );
	OR2X2 OR2X2_63 ( .A(concatenador_counter_2d_0_bF_buf2), .B(micro_hash_synth_2_W_30__1_), .Y(_3528_) );
	INVX1 INVX1_1194 ( .A(micro_hash_synth_2_W_31__1_), .Y(_3529_) );
	NAND2X1 NAND2X1_691 ( .A(concatenador_counter_2d_0_bF_buf1), .B(_3529_), .Y(_3530_) );
	NAND3X1 NAND3X1_222 ( .A(_3439__bF_buf2), .B(_3528_), .C(_3530_), .Y(_3531_) );
	AOI21X1 AOI21X1_886 ( .A(_3527_), .B(_3531_), .C(_3523_), .Y(_3532_) );
	INVX1 INVX1_1195 ( .A(micro_hash_synth_2_W_24__1_), .Y(_3533_) );
	NAND2X1 NAND2X1_692 ( .A(concatenador_counter_2d_0_bF_buf0), .B(micro_hash_synth_2_W_25__1_), .Y(_3534_) );
	OAI21X1 OAI21X1_1263 ( .A(_3533_), .B(concatenador_counter_2d_0_bF_buf12), .C(_3534_), .Y(_3535_) );
	NAND2X1 NAND2X1_693 ( .A(_3440__bF_buf0), .B(_3535_), .Y(_3536_) );
	NAND2X1 NAND2X1_694 ( .A(concatenador_counter_2d_0_bF_buf11), .B(micro_hash_synth_2_W_27__1_), .Y(_3537_) );
	OAI21X1 OAI21X1_1264 ( .A(_4743_), .B(concatenador_counter_2d_0_bF_buf10), .C(_3537_), .Y(_3538_) );
	NAND2X1 NAND2X1_695 ( .A(_3442__bF_buf3), .B(_3538_), .Y(_3539_) );
	NAND3X1 NAND3X1_223 ( .A(_3489__bF_buf3), .B(_3536_), .C(_3539_), .Y(_3540_) );
	OAI21X1 OAI21X1_1265 ( .A(_3540_), .B(_3532_), .C(_3460_), .Y(_3541_) );
	NOR2X1 NOR2X1_566 ( .A(micro_hash_synth_2_W_13__1_), .B(_4733__bF_buf2), .Y(_3542_) );
	OAI21X1 OAI21X1_1266 ( .A(concatenador_counter_2d_0_bF_buf9), .B(micro_hash_synth_2_W_12__1_), .C(concatenador_counter_2d_1_bF_buf6), .Y(_3543_) );
	MUX2X1 MUX2X1_47 ( .A(micro_hash_synth_2_W_15__1_), .B(micro_hash_synth_2_W_14__1_), .S(concatenador_counter_2d_0_bF_buf8), .Y(_3544_) );
	OAI22X1 OAI22X1_516 ( .A(_3544_), .B(concatenador_counter_2d_1_bF_buf5), .C(_3542_), .D(_3543_), .Y(_3545_) );
	INVX1 INVX1_1196 ( .A(micro_hash_synth_2_W_10__1_), .Y(_3546_) );
	NAND2X1 NAND2X1_696 ( .A(concatenador_counter_2d_0_bF_buf7), .B(micro_hash_synth_2_W_11__1_), .Y(_3547_) );
	OAI21X1 OAI21X1_1267 ( .A(_3546_), .B(concatenador_counter_2d_0_bF_buf6), .C(_3547_), .Y(_3548_) );
	NAND2X1 NAND2X1_697 ( .A(_3442__bF_buf2), .B(_3548_), .Y(_3549_) );
	NAND2X1 NAND2X1_698 ( .A(concatenador_counter_2d_0_bF_buf5), .B(micro_hash_synth_2_W_9__1_), .Y(_3550_) );
	OAI21X1 OAI21X1_1268 ( .A(_4802_), .B(concatenador_counter_2d_0_bF_buf4), .C(_3550_), .Y(_3551_) );
	NAND2X1 NAND2X1_699 ( .A(_3440__bF_buf4), .B(_3551_), .Y(_3552_) );
	NAND3X1 NAND3X1_224 ( .A(_3489__bF_buf2), .B(_3549_), .C(_3552_), .Y(_3553_) );
	AOI21X1 AOI21X1_887 ( .A(_3443__bF_buf0), .B(_3545_), .C(_3553_), .Y(_3554_) );
	INVX1 INVX1_1197 ( .A(micro_hash_synth_2_W_5__1_), .Y(_3555_) );
	NAND2X1 NAND2X1_700 ( .A(concatenador_counter_2d_0_bF_buf3), .B(_3555_), .Y(_3556_) );
	OR2X2 OR2X2_64 ( .A(concatenador_counter_2d_0_bF_buf2), .B(micro_hash_synth_2_W_4__1_), .Y(_3557_) );
	NAND3X1 NAND3X1_225 ( .A(concatenador_counter_2d_1_bF_buf4), .B(_3557_), .C(_3556_), .Y(_3558_) );
	OR2X2 OR2X2_65 ( .A(concatenador_counter_2d_0_bF_buf1), .B(micro_hash_synth_2_W_6__1_), .Y(_3559_) );
	INVX1 INVX1_1198 ( .A(micro_hash_synth_2_W_7__1_), .Y(_3560_) );
	NAND2X1 NAND2X1_701 ( .A(concatenador_counter_2d_0_bF_buf0), .B(_3560_), .Y(_3561_) );
	NAND3X1 NAND3X1_226 ( .A(_3439__bF_buf1), .B(_3559_), .C(_3561_), .Y(_3562_) );
	AOI21X1 AOI21X1_888 ( .A(_3558_), .B(_3562_), .C(_3523_), .Y(_3563_) );
	NAND2X1 NAND2X1_702 ( .A(concatenador_counter_2d_0_bF_buf12), .B(micro_hash_synth_2_W_1__1_), .Y(_3564_) );
	OAI21X1 OAI21X1_1269 ( .A(_4842_), .B(concatenador_counter_2d_0_bF_buf11), .C(_3564_), .Y(_3565_) );
	NAND2X1 NAND2X1_703 ( .A(_3440__bF_buf3), .B(_3565_), .Y(_3566_) );
	NAND2X1 NAND2X1_704 ( .A(concatenador_counter_2d_0_bF_buf10), .B(micro_hash_synth_2_W_3__1_), .Y(_3567_) );
	OAI21X1 OAI21X1_1270 ( .A(_4850_), .B(concatenador_counter_2d_0_bF_buf9), .C(_3567_), .Y(_3568_) );
	NAND2X1 NAND2X1_705 ( .A(_3442__bF_buf1), .B(_3568_), .Y(_3569_) );
	NAND3X1 NAND3X1_227 ( .A(_3453__bF_buf0), .B(_3566_), .C(_3569_), .Y(_3570_) );
	OAI21X1 OAI21X1_1271 ( .A(_3570_), .B(_3563_), .C(_3490_), .Y(_3571_) );
	OAI22X1 OAI22X1_517 ( .A(_3541_), .B(_3522_), .C(_3554_), .D(_3571_), .Y(_3572_) );
	AND2X2 AND2X2_99 ( .A(micro_hash_synth_2_k_1_), .B(micro_hash_synth_2_x_1_), .Y(_3573_) );
	NOR2X1 NOR2X1_567 ( .A(micro_hash_synth_2_k_1_), .B(micro_hash_synth_2_x_1_), .Y(_3574_) );
	NOR2X1 NOR2X1_568 ( .A(_3574_), .B(_3573_), .Y(_3575_) );
	NAND2X1 NAND2X1_706 ( .A(_3575_), .B(_3572_), .Y(_3576_) );
	NAND2X1 NAND2X1_707 ( .A(_3443__bF_buf5), .B(_3512_), .Y(_3577_) );
	AOI21X1 AOI21X1_889 ( .A(_3440__bF_buf2), .B(_3519_), .C(_3489__bF_buf1), .Y(_3578_) );
	NAND3X1 NAND3X1_228 ( .A(_3516_), .B(_3578_), .C(_3577_), .Y(_3579_) );
	NOR2X1 NOR2X1_569 ( .A(micro_hash_synth_2_W_29__1_), .B(_4733__bF_buf1), .Y(_3580_) );
	OAI21X1 OAI21X1_1272 ( .A(concatenador_counter_2d_0_bF_buf8), .B(micro_hash_synth_2_W_28__1_), .C(concatenador_counter_2d_1_bF_buf3), .Y(_3581_) );
	MUX2X1 MUX2X1_48 ( .A(micro_hash_synth_2_W_31__1_), .B(micro_hash_synth_2_W_30__1_), .S(concatenador_counter_2d_0_bF_buf7), .Y(_3582_) );
endmodule
